module DRAM (
input wire [15:0] address,
input clock,
input wire [7:0] data,
input wren,
output reg [7:0] q);
reg [7:0] DRAM[524287:0];

initial begin
DRAM[0] = 8'b1011000;
DRAM[1] = 8'b1011000;
DRAM[2] = 8'b1011001;
DRAM[3] = 8'b1011001;
DRAM[4] = 8'b1011010;
DRAM[5] = 8'b1011011;
DRAM[6] = 8'b1011100;
DRAM[7] = 8'b1011100;
DRAM[8] = 8'b1011100;
DRAM[9] = 8'b1011011;
DRAM[10] = 8'b1011011;
DRAM[11] = 8'b1011100;
DRAM[12] = 8'b1011111;
DRAM[13] = 8'b1100001;
DRAM[14] = 8'b1100001;
DRAM[15] = 8'b1100000;
DRAM[16] = 8'b1011111;
DRAM[17] = 8'b1100000;
DRAM[18] = 8'b1100010;
DRAM[19] = 8'b1100011;
DRAM[20] = 8'b1100100;
DRAM[21] = 8'b1100011;
DRAM[22] = 8'b1100010;
DRAM[23] = 8'b1100001;
DRAM[24] = 8'b1100101;
DRAM[25] = 8'b1100101;
DRAM[26] = 8'b1100101;
DRAM[27] = 8'b1100110;
DRAM[28] = 8'b1100110;
DRAM[29] = 8'b1100111;
DRAM[30] = 8'b1100111;
DRAM[31] = 8'b1100111;
DRAM[32] = 8'b1100110;
DRAM[33] = 8'b1100110;
DRAM[34] = 8'b1100111;
DRAM[35] = 8'b1100111;
DRAM[36] = 8'b1100111;
DRAM[37] = 8'b1100111;
DRAM[38] = 8'b1100111;
DRAM[39] = 8'b1101000;
DRAM[40] = 8'b1101011;
DRAM[41] = 8'b1101011;
DRAM[42] = 8'b1101011;
DRAM[43] = 8'b1101011;
DRAM[44] = 8'b1101011;
DRAM[45] = 8'b1101011;
DRAM[46] = 8'b1101011;
DRAM[47] = 8'b1101011;
DRAM[48] = 8'b1101100;
DRAM[49] = 8'b1101100;
DRAM[50] = 8'b1101100;
DRAM[51] = 8'b1101100;
DRAM[52] = 8'b1101100;
DRAM[53] = 8'b1101100;
DRAM[54] = 8'b1101100;
DRAM[55] = 8'b1101100;
DRAM[56] = 8'b1101101;
DRAM[57] = 8'b1101101;
DRAM[58] = 8'b1101101;
DRAM[59] = 8'b1101101;
DRAM[60] = 8'b1101101;
DRAM[61] = 8'b1101101;
DRAM[62] = 8'b1101101;
DRAM[63] = 8'b1101101;
DRAM[64] = 8'b1101110;
DRAM[65] = 8'b1101110;
DRAM[66] = 8'b1101110;
DRAM[67] = 8'b1101101;
DRAM[68] = 8'b1101101;
DRAM[69] = 8'b1101100;
DRAM[70] = 8'b1101100;
DRAM[71] = 8'b1101011;
DRAM[72] = 8'b1101100;
DRAM[73] = 8'b1101100;
DRAM[74] = 8'b1101101;
DRAM[75] = 8'b1101101;
DRAM[76] = 8'b1101101;
DRAM[77] = 8'b1101100;
DRAM[78] = 8'b1101011;
DRAM[79] = 8'b1101010;
DRAM[80] = 8'b1101100;
DRAM[81] = 8'b1101011;
DRAM[82] = 8'b1101010;
DRAM[83] = 8'b1101001;
DRAM[84] = 8'b1101001;
DRAM[85] = 8'b1101001;
DRAM[86] = 8'b1101001;
DRAM[87] = 8'b1101010;
DRAM[88] = 8'b1101010;
DRAM[89] = 8'b1101010;
DRAM[90] = 8'b1101010;
DRAM[91] = 8'b1101010;
DRAM[92] = 8'b1101010;
DRAM[93] = 8'b1101010;
DRAM[94] = 8'b1101010;
DRAM[95] = 8'b1101010;
DRAM[96] = 8'b1101101;
DRAM[97] = 8'b1101101;
DRAM[98] = 8'b1101100;
DRAM[99] = 8'b1101100;
DRAM[100] = 8'b1101100;
DRAM[101] = 8'b1101101;
DRAM[102] = 8'b1101110;
DRAM[103] = 8'b1101111;
DRAM[104] = 8'b1101011;
DRAM[105] = 8'b1101011;
DRAM[106] = 8'b1101010;
DRAM[107] = 8'b1101010;
DRAM[108] = 8'b1101010;
DRAM[109] = 8'b1101001;
DRAM[110] = 8'b1101001;
DRAM[111] = 8'b1101001;
DRAM[112] = 8'b1101001;
DRAM[113] = 8'b1101001;
DRAM[114] = 8'b1101001;
DRAM[115] = 8'b1101001;
DRAM[116] = 8'b1101001;
DRAM[117] = 8'b1101001;
DRAM[118] = 8'b1101001;
DRAM[119] = 8'b1101001;
DRAM[120] = 8'b1101000;
DRAM[121] = 8'b1101000;
DRAM[122] = 8'b1101000;
DRAM[123] = 8'b1101000;
DRAM[124] = 8'b1101000;
DRAM[125] = 8'b1101000;
DRAM[126] = 8'b1101000;
DRAM[127] = 8'b1101000;
DRAM[128] = 8'b1100111;
DRAM[129] = 8'b1101000;
DRAM[130] = 8'b1101000;
DRAM[131] = 8'b1101001;
DRAM[132] = 8'b1101001;
DRAM[133] = 8'b1101010;
DRAM[134] = 8'b1101010;
DRAM[135] = 8'b1101010;
DRAM[136] = 8'b1100111;
DRAM[137] = 8'b1101000;
DRAM[138] = 8'b1101001;
DRAM[139] = 8'b1101010;
DRAM[140] = 8'b1101010;
DRAM[141] = 8'b1101010;
DRAM[142] = 8'b1101001;
DRAM[143] = 8'b1101001;
DRAM[144] = 8'b1101001;
DRAM[145] = 8'b1101010;
DRAM[146] = 8'b1101010;
DRAM[147] = 8'b1101011;
DRAM[148] = 8'b1101011;
DRAM[149] = 8'b1101010;
DRAM[150] = 8'b1101010;
DRAM[151] = 8'b1101001;
DRAM[152] = 8'b1101000;
DRAM[153] = 8'b1101000;
DRAM[154] = 8'b1101000;
DRAM[155] = 8'b1101000;
DRAM[156] = 8'b1101000;
DRAM[157] = 8'b1101000;
DRAM[158] = 8'b1101000;
DRAM[159] = 8'b1101000;
DRAM[160] = 8'b1100110;
DRAM[161] = 8'b1100110;
DRAM[162] = 8'b1100110;
DRAM[163] = 8'b1100110;
DRAM[164] = 8'b1100101;
DRAM[165] = 8'b1100100;
DRAM[166] = 8'b1100011;
DRAM[167] = 8'b1100010;
DRAM[168] = 8'b1100100;
DRAM[169] = 8'b1100010;
DRAM[170] = 8'b1100001;
DRAM[171] = 8'b1100000;
DRAM[172] = 8'b1011111;
DRAM[173] = 8'b1100000;
DRAM[174] = 8'b1100001;
DRAM[175] = 8'b1100001;
DRAM[176] = 8'b1011111;
DRAM[177] = 8'b1011111;
DRAM[178] = 8'b1011110;
DRAM[179] = 8'b1011110;
DRAM[180] = 8'b1011110;
DRAM[181] = 8'b1011101;
DRAM[182] = 8'b1011101;
DRAM[183] = 8'b1011101;
DRAM[184] = 8'b1011011;
DRAM[185] = 8'b1011011;
DRAM[186] = 8'b1011010;
DRAM[187] = 8'b1011001;
DRAM[188] = 8'b1011000;
DRAM[189] = 8'b1011000;
DRAM[190] = 8'b1010111;
DRAM[191] = 8'b1010111;
DRAM[192] = 8'b1010101;
DRAM[193] = 8'b1010101;
DRAM[194] = 8'b1010101;
DRAM[195] = 8'b1010101;
DRAM[196] = 8'b1010101;
DRAM[197] = 8'b1010101;
DRAM[198] = 8'b1010101;
DRAM[199] = 8'b1010101;
DRAM[200] = 8'b1010011;
DRAM[201] = 8'b1010011;
DRAM[202] = 8'b1010010;
DRAM[203] = 8'b1010010;
DRAM[204] = 8'b1010010;
DRAM[205] = 8'b1010001;
DRAM[206] = 8'b1010001;
DRAM[207] = 8'b1010001;
DRAM[208] = 8'b1010000;
DRAM[209] = 8'b1010000;
DRAM[210] = 8'b1010000;
DRAM[211] = 8'b1001111;
DRAM[212] = 8'b1001111;
DRAM[213] = 8'b1001110;
DRAM[214] = 8'b1001110;
DRAM[215] = 8'b1001110;
DRAM[216] = 8'b1001001;
DRAM[217] = 8'b1001010;
DRAM[218] = 8'b1001010;
DRAM[219] = 8'b1001011;
DRAM[220] = 8'b1001011;
DRAM[221] = 8'b1001010;
DRAM[222] = 8'b1001001;
DRAM[223] = 8'b1001000;
DRAM[224] = 8'b1000111;
DRAM[225] = 8'b1000111;
DRAM[226] = 8'b1000110;
DRAM[227] = 8'b1000110;
DRAM[228] = 8'b1000110;
DRAM[229] = 8'b1000101;
DRAM[230] = 8'b1000101;
DRAM[231] = 8'b1000101;
DRAM[232] = 8'b1000100;
DRAM[233] = 8'b1000100;
DRAM[234] = 8'b1000100;
DRAM[235] = 8'b1000011;
DRAM[236] = 8'b1000011;
DRAM[237] = 8'b1000010;
DRAM[238] = 8'b1000010;
DRAM[239] = 8'b1000010;
DRAM[240] = 8'b1000010;
DRAM[241] = 8'b1000010;
DRAM[242] = 8'b1000010;
DRAM[243] = 8'b1000001;
DRAM[244] = 8'b1000001;
DRAM[245] = 8'b1000000;
DRAM[246] = 8'b1000000;
DRAM[247] = 8'b1000000;
DRAM[248] = 8'b1000000;
DRAM[249] = 8'b1000000;
DRAM[250] = 8'b1000000;
DRAM[251] = 8'b111111;
DRAM[252] = 8'b111111;
DRAM[253] = 8'b111111;
DRAM[254] = 8'b111110;
DRAM[255] = 8'b111110;
DRAM[256] = 8'b1011000;
DRAM[257] = 8'b1011000;
DRAM[258] = 8'b1011001;
DRAM[259] = 8'b1011010;
DRAM[260] = 8'b1011011;
DRAM[261] = 8'b1011011;
DRAM[262] = 8'b1011100;
DRAM[263] = 8'b1011100;
DRAM[264] = 8'b1011100;
DRAM[265] = 8'b1011011;
DRAM[266] = 8'b1011011;
DRAM[267] = 8'b1011101;
DRAM[268] = 8'b1100000;
DRAM[269] = 8'b1100001;
DRAM[270] = 8'b1100001;
DRAM[271] = 8'b1100000;
DRAM[272] = 8'b1100001;
DRAM[273] = 8'b1100001;
DRAM[274] = 8'b1100010;
DRAM[275] = 8'b1100011;
DRAM[276] = 8'b1100011;
DRAM[277] = 8'b1100011;
DRAM[278] = 8'b1100011;
DRAM[279] = 8'b1100011;
DRAM[280] = 8'b1100100;
DRAM[281] = 8'b1100100;
DRAM[282] = 8'b1100100;
DRAM[283] = 8'b1100101;
DRAM[284] = 8'b1100101;
DRAM[285] = 8'b1100101;
DRAM[286] = 8'b1100110;
DRAM[287] = 8'b1100110;
DRAM[288] = 8'b1100110;
DRAM[289] = 8'b1100111;
DRAM[290] = 8'b1100111;
DRAM[291] = 8'b1100111;
DRAM[292] = 8'b1100111;
DRAM[293] = 8'b1101000;
DRAM[294] = 8'b1101000;
DRAM[295] = 8'b1101000;
DRAM[296] = 8'b1101011;
DRAM[297] = 8'b1101011;
DRAM[298] = 8'b1101011;
DRAM[299] = 8'b1101011;
DRAM[300] = 8'b1101011;
DRAM[301] = 8'b1101011;
DRAM[302] = 8'b1101011;
DRAM[303] = 8'b1101011;
DRAM[304] = 8'b1101100;
DRAM[305] = 8'b1101100;
DRAM[306] = 8'b1101100;
DRAM[307] = 8'b1101100;
DRAM[308] = 8'b1101100;
DRAM[309] = 8'b1101100;
DRAM[310] = 8'b1101100;
DRAM[311] = 8'b1101100;
DRAM[312] = 8'b1101101;
DRAM[313] = 8'b1101101;
DRAM[314] = 8'b1101101;
DRAM[315] = 8'b1101101;
DRAM[316] = 8'b1101101;
DRAM[317] = 8'b1101101;
DRAM[318] = 8'b1101101;
DRAM[319] = 8'b1101101;
DRAM[320] = 8'b1101110;
DRAM[321] = 8'b1101110;
DRAM[322] = 8'b1101110;
DRAM[323] = 8'b1101101;
DRAM[324] = 8'b1101101;
DRAM[325] = 8'b1101101;
DRAM[326] = 8'b1101100;
DRAM[327] = 8'b1101100;
DRAM[328] = 8'b1101100;
DRAM[329] = 8'b1101101;
DRAM[330] = 8'b1101101;
DRAM[331] = 8'b1101101;
DRAM[332] = 8'b1101101;
DRAM[333] = 8'b1101100;
DRAM[334] = 8'b1101011;
DRAM[335] = 8'b1101010;
DRAM[336] = 8'b1101100;
DRAM[337] = 8'b1101011;
DRAM[338] = 8'b1101011;
DRAM[339] = 8'b1101010;
DRAM[340] = 8'b1101001;
DRAM[341] = 8'b1101001;
DRAM[342] = 8'b1101010;
DRAM[343] = 8'b1101010;
DRAM[344] = 8'b1101010;
DRAM[345] = 8'b1101010;
DRAM[346] = 8'b1101010;
DRAM[347] = 8'b1101010;
DRAM[348] = 8'b1101010;
DRAM[349] = 8'b1101010;
DRAM[350] = 8'b1101010;
DRAM[351] = 8'b1101010;
DRAM[352] = 8'b1101100;
DRAM[353] = 8'b1101100;
DRAM[354] = 8'b1101100;
DRAM[355] = 8'b1101100;
DRAM[356] = 8'b1101100;
DRAM[357] = 8'b1101101;
DRAM[358] = 8'b1101110;
DRAM[359] = 8'b1101110;
DRAM[360] = 8'b1101011;
DRAM[361] = 8'b1101011;
DRAM[362] = 8'b1101011;
DRAM[363] = 8'b1101010;
DRAM[364] = 8'b1101010;
DRAM[365] = 8'b1101010;
DRAM[366] = 8'b1101001;
DRAM[367] = 8'b1101001;
DRAM[368] = 8'b1101001;
DRAM[369] = 8'b1101001;
DRAM[370] = 8'b1101001;
DRAM[371] = 8'b1101001;
DRAM[372] = 8'b1101001;
DRAM[373] = 8'b1101001;
DRAM[374] = 8'b1101001;
DRAM[375] = 8'b1101001;
DRAM[376] = 8'b1101000;
DRAM[377] = 8'b1101000;
DRAM[378] = 8'b1101000;
DRAM[379] = 8'b1101000;
DRAM[380] = 8'b1101000;
DRAM[381] = 8'b1101000;
DRAM[382] = 8'b1101000;
DRAM[383] = 8'b1101000;
DRAM[384] = 8'b1101000;
DRAM[385] = 8'b1101000;
DRAM[386] = 8'b1101001;
DRAM[387] = 8'b1101001;
DRAM[388] = 8'b1101001;
DRAM[389] = 8'b1101010;
DRAM[390] = 8'b1101010;
DRAM[391] = 8'b1101010;
DRAM[392] = 8'b1100111;
DRAM[393] = 8'b1101000;
DRAM[394] = 8'b1101001;
DRAM[395] = 8'b1101010;
DRAM[396] = 8'b1101010;
DRAM[397] = 8'b1101010;
DRAM[398] = 8'b1101010;
DRAM[399] = 8'b1101001;
DRAM[400] = 8'b1101000;
DRAM[401] = 8'b1101000;
DRAM[402] = 8'b1101001;
DRAM[403] = 8'b1101001;
DRAM[404] = 8'b1101001;
DRAM[405] = 8'b1101001;
DRAM[406] = 8'b1101000;
DRAM[407] = 8'b1101000;
DRAM[408] = 8'b1100111;
DRAM[409] = 8'b1100111;
DRAM[410] = 8'b1100111;
DRAM[411] = 8'b1100111;
DRAM[412] = 8'b1100111;
DRAM[413] = 8'b1100111;
DRAM[414] = 8'b1100111;
DRAM[415] = 8'b1100111;
DRAM[416] = 8'b1100111;
DRAM[417] = 8'b1100111;
DRAM[418] = 8'b1100111;
DRAM[419] = 8'b1100110;
DRAM[420] = 8'b1100110;
DRAM[421] = 8'b1100100;
DRAM[422] = 8'b1100011;
DRAM[423] = 8'b1100010;
DRAM[424] = 8'b1100100;
DRAM[425] = 8'b1100011;
DRAM[426] = 8'b1100001;
DRAM[427] = 8'b1100000;
DRAM[428] = 8'b1100000;
DRAM[429] = 8'b1100000;
DRAM[430] = 8'b1100001;
DRAM[431] = 8'b1100010;
DRAM[432] = 8'b1011111;
DRAM[433] = 8'b1011111;
DRAM[434] = 8'b1011111;
DRAM[435] = 8'b1011110;
DRAM[436] = 8'b1011110;
DRAM[437] = 8'b1011110;
DRAM[438] = 8'b1011101;
DRAM[439] = 8'b1011101;
DRAM[440] = 8'b1011011;
DRAM[441] = 8'b1011011;
DRAM[442] = 8'b1011011;
DRAM[443] = 8'b1011010;
DRAM[444] = 8'b1011001;
DRAM[445] = 8'b1011000;
DRAM[446] = 8'b1011000;
DRAM[447] = 8'b1010111;
DRAM[448] = 8'b1010101;
DRAM[449] = 8'b1010101;
DRAM[450] = 8'b1010101;
DRAM[451] = 8'b1010101;
DRAM[452] = 8'b1010101;
DRAM[453] = 8'b1010101;
DRAM[454] = 8'b1010101;
DRAM[455] = 8'b1010101;
DRAM[456] = 8'b1010011;
DRAM[457] = 8'b1010011;
DRAM[458] = 8'b1010011;
DRAM[459] = 8'b1010010;
DRAM[460] = 8'b1010010;
DRAM[461] = 8'b1010010;
DRAM[462] = 8'b1010001;
DRAM[463] = 8'b1010001;
DRAM[464] = 8'b1010000;
DRAM[465] = 8'b1010000;
DRAM[466] = 8'b1010000;
DRAM[467] = 8'b1001111;
DRAM[468] = 8'b1001111;
DRAM[469] = 8'b1001111;
DRAM[470] = 8'b1001110;
DRAM[471] = 8'b1001110;
DRAM[472] = 8'b1001011;
DRAM[473] = 8'b1001100;
DRAM[474] = 8'b1001100;
DRAM[475] = 8'b1001100;
DRAM[476] = 8'b1001011;
DRAM[477] = 8'b1001010;
DRAM[478] = 8'b1001001;
DRAM[479] = 8'b1001001;
DRAM[480] = 8'b1000111;
DRAM[481] = 8'b1000111;
DRAM[482] = 8'b1000111;
DRAM[483] = 8'b1000110;
DRAM[484] = 8'b1000110;
DRAM[485] = 8'b1000110;
DRAM[486] = 8'b1000101;
DRAM[487] = 8'b1000101;
DRAM[488] = 8'b1000101;
DRAM[489] = 8'b1000101;
DRAM[490] = 8'b1000101;
DRAM[491] = 8'b1000101;
DRAM[492] = 8'b1000100;
DRAM[493] = 8'b1000100;
DRAM[494] = 8'b1000011;
DRAM[495] = 8'b1000011;
DRAM[496] = 8'b1000010;
DRAM[497] = 8'b1000010;
DRAM[498] = 8'b1000010;
DRAM[499] = 8'b1000001;
DRAM[500] = 8'b1000001;
DRAM[501] = 8'b1000001;
DRAM[502] = 8'b1000000;
DRAM[503] = 8'b1000000;
DRAM[504] = 8'b1000000;
DRAM[505] = 8'b111111;
DRAM[506] = 8'b111111;
DRAM[507] = 8'b111111;
DRAM[508] = 8'b111110;
DRAM[509] = 8'b111110;
DRAM[510] = 8'b111110;
DRAM[511] = 8'b111110;
DRAM[512] = 8'b1011001;
DRAM[513] = 8'b1011001;
DRAM[514] = 8'b1011010;
DRAM[515] = 8'b1011010;
DRAM[516] = 8'b1011011;
DRAM[517] = 8'b1011100;
DRAM[518] = 8'b1011101;
DRAM[519] = 8'b1011101;
DRAM[520] = 8'b1011101;
DRAM[521] = 8'b1011100;
DRAM[522] = 8'b1011100;
DRAM[523] = 8'b1011101;
DRAM[524] = 8'b1100000;
DRAM[525] = 8'b1100010;
DRAM[526] = 8'b1100010;
DRAM[527] = 8'b1100001;
DRAM[528] = 8'b1100011;
DRAM[529] = 8'b1100011;
DRAM[530] = 8'b1100010;
DRAM[531] = 8'b1100010;
DRAM[532] = 8'b1100011;
DRAM[533] = 8'b1100100;
DRAM[534] = 8'b1100100;
DRAM[535] = 8'b1100101;
DRAM[536] = 8'b1100011;
DRAM[537] = 8'b1100011;
DRAM[538] = 8'b1100100;
DRAM[539] = 8'b1100100;
DRAM[540] = 8'b1100100;
DRAM[541] = 8'b1100101;
DRAM[542] = 8'b1100101;
DRAM[543] = 8'b1100101;
DRAM[544] = 8'b1100111;
DRAM[545] = 8'b1100111;
DRAM[546] = 8'b1100111;
DRAM[547] = 8'b1101000;
DRAM[548] = 8'b1101000;
DRAM[549] = 8'b1101001;
DRAM[550] = 8'b1101001;
DRAM[551] = 8'b1101001;
DRAM[552] = 8'b1101100;
DRAM[553] = 8'b1101100;
DRAM[554] = 8'b1101100;
DRAM[555] = 8'b1101100;
DRAM[556] = 8'b1101100;
DRAM[557] = 8'b1101100;
DRAM[558] = 8'b1101100;
DRAM[559] = 8'b1101100;
DRAM[560] = 8'b1101101;
DRAM[561] = 8'b1101101;
DRAM[562] = 8'b1101101;
DRAM[563] = 8'b1101101;
DRAM[564] = 8'b1101101;
DRAM[565] = 8'b1101101;
DRAM[566] = 8'b1101101;
DRAM[567] = 8'b1101101;
DRAM[568] = 8'b1101110;
DRAM[569] = 8'b1101110;
DRAM[570] = 8'b1101110;
DRAM[571] = 8'b1101110;
DRAM[572] = 8'b1101110;
DRAM[573] = 8'b1101110;
DRAM[574] = 8'b1101110;
DRAM[575] = 8'b1101110;
DRAM[576] = 8'b1101111;
DRAM[577] = 8'b1101111;
DRAM[578] = 8'b1101110;
DRAM[579] = 8'b1101110;
DRAM[580] = 8'b1101110;
DRAM[581] = 8'b1101101;
DRAM[582] = 8'b1101101;
DRAM[583] = 8'b1101101;
DRAM[584] = 8'b1101101;
DRAM[585] = 8'b1101101;
DRAM[586] = 8'b1101110;
DRAM[587] = 8'b1101110;
DRAM[588] = 8'b1101101;
DRAM[589] = 8'b1101101;
DRAM[590] = 8'b1101100;
DRAM[591] = 8'b1101011;
DRAM[592] = 8'b1101101;
DRAM[593] = 8'b1101100;
DRAM[594] = 8'b1101011;
DRAM[595] = 8'b1101010;
DRAM[596] = 8'b1101010;
DRAM[597] = 8'b1101010;
DRAM[598] = 8'b1101010;
DRAM[599] = 8'b1101011;
DRAM[600] = 8'b1101011;
DRAM[601] = 8'b1101011;
DRAM[602] = 8'b1101011;
DRAM[603] = 8'b1101011;
DRAM[604] = 8'b1101011;
DRAM[605] = 8'b1101011;
DRAM[606] = 8'b1101011;
DRAM[607] = 8'b1101011;
DRAM[608] = 8'b1101100;
DRAM[609] = 8'b1101011;
DRAM[610] = 8'b1101011;
DRAM[611] = 8'b1101011;
DRAM[612] = 8'b1101011;
DRAM[613] = 8'b1101100;
DRAM[614] = 8'b1101101;
DRAM[615] = 8'b1101110;
DRAM[616] = 8'b1101100;
DRAM[617] = 8'b1101100;
DRAM[618] = 8'b1101011;
DRAM[619] = 8'b1101011;
DRAM[620] = 8'b1101011;
DRAM[621] = 8'b1101010;
DRAM[622] = 8'b1101010;
DRAM[623] = 8'b1101010;
DRAM[624] = 8'b1101010;
DRAM[625] = 8'b1101010;
DRAM[626] = 8'b1101010;
DRAM[627] = 8'b1101010;
DRAM[628] = 8'b1101010;
DRAM[629] = 8'b1101010;
DRAM[630] = 8'b1101010;
DRAM[631] = 8'b1101010;
DRAM[632] = 8'b1101001;
DRAM[633] = 8'b1101001;
DRAM[634] = 8'b1101001;
DRAM[635] = 8'b1101001;
DRAM[636] = 8'b1101001;
DRAM[637] = 8'b1101001;
DRAM[638] = 8'b1101001;
DRAM[639] = 8'b1101001;
DRAM[640] = 8'b1101001;
DRAM[641] = 8'b1101001;
DRAM[642] = 8'b1101001;
DRAM[643] = 8'b1101010;
DRAM[644] = 8'b1101010;
DRAM[645] = 8'b1101010;
DRAM[646] = 8'b1101011;
DRAM[647] = 8'b1101011;
DRAM[648] = 8'b1101000;
DRAM[649] = 8'b1101001;
DRAM[650] = 8'b1101010;
DRAM[651] = 8'b1101010;
DRAM[652] = 8'b1101011;
DRAM[653] = 8'b1101011;
DRAM[654] = 8'b1101010;
DRAM[655] = 8'b1101010;
DRAM[656] = 8'b1100111;
DRAM[657] = 8'b1100111;
DRAM[658] = 8'b1101000;
DRAM[659] = 8'b1101000;
DRAM[660] = 8'b1101000;
DRAM[661] = 8'b1101000;
DRAM[662] = 8'b1100111;
DRAM[663] = 8'b1100111;
DRAM[664] = 8'b1100110;
DRAM[665] = 8'b1100110;
DRAM[666] = 8'b1100110;
DRAM[667] = 8'b1100110;
DRAM[668] = 8'b1100110;
DRAM[669] = 8'b1100110;
DRAM[670] = 8'b1100110;
DRAM[671] = 8'b1100110;
DRAM[672] = 8'b1100111;
DRAM[673] = 8'b1100111;
DRAM[674] = 8'b1100111;
DRAM[675] = 8'b1100111;
DRAM[676] = 8'b1100110;
DRAM[677] = 8'b1100101;
DRAM[678] = 8'b1100100;
DRAM[679] = 8'b1100011;
DRAM[680] = 8'b1100100;
DRAM[681] = 8'b1100011;
DRAM[682] = 8'b1100010;
DRAM[683] = 8'b1100001;
DRAM[684] = 8'b1100001;
DRAM[685] = 8'b1100001;
DRAM[686] = 8'b1100001;
DRAM[687] = 8'b1100010;
DRAM[688] = 8'b1100000;
DRAM[689] = 8'b1100000;
DRAM[690] = 8'b1011111;
DRAM[691] = 8'b1011111;
DRAM[692] = 8'b1011111;
DRAM[693] = 8'b1011110;
DRAM[694] = 8'b1011110;
DRAM[695] = 8'b1011110;
DRAM[696] = 8'b1011100;
DRAM[697] = 8'b1011100;
DRAM[698] = 8'b1011011;
DRAM[699] = 8'b1011011;
DRAM[700] = 8'b1011010;
DRAM[701] = 8'b1011001;
DRAM[702] = 8'b1011000;
DRAM[703] = 8'b1011000;
DRAM[704] = 8'b1010110;
DRAM[705] = 8'b1010110;
DRAM[706] = 8'b1010110;
DRAM[707] = 8'b1010110;
DRAM[708] = 8'b1010110;
DRAM[709] = 8'b1010110;
DRAM[710] = 8'b1010110;
DRAM[711] = 8'b1010110;
DRAM[712] = 8'b1010100;
DRAM[713] = 8'b1010100;
DRAM[714] = 8'b1010011;
DRAM[715] = 8'b1010011;
DRAM[716] = 8'b1010011;
DRAM[717] = 8'b1010010;
DRAM[718] = 8'b1010010;
DRAM[719] = 8'b1010010;
DRAM[720] = 8'b1010000;
DRAM[721] = 8'b1010000;
DRAM[722] = 8'b1010000;
DRAM[723] = 8'b1010000;
DRAM[724] = 8'b1001111;
DRAM[725] = 8'b1001111;
DRAM[726] = 8'b1001111;
DRAM[727] = 8'b1001110;
DRAM[728] = 8'b1001110;
DRAM[729] = 8'b1001110;
DRAM[730] = 8'b1001110;
DRAM[731] = 8'b1001110;
DRAM[732] = 8'b1001101;
DRAM[733] = 8'b1001011;
DRAM[734] = 8'b1001010;
DRAM[735] = 8'b1001001;
DRAM[736] = 8'b1001000;
DRAM[737] = 8'b1001000;
DRAM[738] = 8'b1000111;
DRAM[739] = 8'b1000111;
DRAM[740] = 8'b1000111;
DRAM[741] = 8'b1000110;
DRAM[742] = 8'b1000110;
DRAM[743] = 8'b1000110;
DRAM[744] = 8'b1000111;
DRAM[745] = 8'b1000111;
DRAM[746] = 8'b1000110;
DRAM[747] = 8'b1000110;
DRAM[748] = 8'b1000101;
DRAM[749] = 8'b1000101;
DRAM[750] = 8'b1000101;
DRAM[751] = 8'b1000101;
DRAM[752] = 8'b1000010;
DRAM[753] = 8'b1000010;
DRAM[754] = 8'b1000010;
DRAM[755] = 8'b1000010;
DRAM[756] = 8'b1000001;
DRAM[757] = 8'b1000001;
DRAM[758] = 8'b1000001;
DRAM[759] = 8'b1000000;
DRAM[760] = 8'b111111;
DRAM[761] = 8'b111111;
DRAM[762] = 8'b111111;
DRAM[763] = 8'b111110;
DRAM[764] = 8'b111110;
DRAM[765] = 8'b111101;
DRAM[766] = 8'b111101;
DRAM[767] = 8'b111101;
DRAM[768] = 8'b1011010;
DRAM[769] = 8'b1011010;
DRAM[770] = 8'b1011010;
DRAM[771] = 8'b1011011;
DRAM[772] = 8'b1011100;
DRAM[773] = 8'b1011101;
DRAM[774] = 8'b1011101;
DRAM[775] = 8'b1011110;
DRAM[776] = 8'b1011110;
DRAM[777] = 8'b1011101;
DRAM[778] = 8'b1011100;
DRAM[779] = 8'b1011110;
DRAM[780] = 8'b1100001;
DRAM[781] = 8'b1100011;
DRAM[782] = 8'b1100011;
DRAM[783] = 8'b1100010;
DRAM[784] = 8'b1100101;
DRAM[785] = 8'b1100100;
DRAM[786] = 8'b1100011;
DRAM[787] = 8'b1100010;
DRAM[788] = 8'b1100011;
DRAM[789] = 8'b1100100;
DRAM[790] = 8'b1100110;
DRAM[791] = 8'b1100111;
DRAM[792] = 8'b1100100;
DRAM[793] = 8'b1100100;
DRAM[794] = 8'b1100101;
DRAM[795] = 8'b1100101;
DRAM[796] = 8'b1100101;
DRAM[797] = 8'b1100110;
DRAM[798] = 8'b1100110;
DRAM[799] = 8'b1100110;
DRAM[800] = 8'b1100111;
DRAM[801] = 8'b1100111;
DRAM[802] = 8'b1101000;
DRAM[803] = 8'b1101000;
DRAM[804] = 8'b1101001;
DRAM[805] = 8'b1101010;
DRAM[806] = 8'b1101010;
DRAM[807] = 8'b1101010;
DRAM[808] = 8'b1101100;
DRAM[809] = 8'b1101100;
DRAM[810] = 8'b1101100;
DRAM[811] = 8'b1101100;
DRAM[812] = 8'b1101101;
DRAM[813] = 8'b1101101;
DRAM[814] = 8'b1101101;
DRAM[815] = 8'b1101101;
DRAM[816] = 8'b1101110;
DRAM[817] = 8'b1101110;
DRAM[818] = 8'b1101110;
DRAM[819] = 8'b1101110;
DRAM[820] = 8'b1101110;
DRAM[821] = 8'b1101110;
DRAM[822] = 8'b1101110;
DRAM[823] = 8'b1101110;
DRAM[824] = 8'b1101111;
DRAM[825] = 8'b1101111;
DRAM[826] = 8'b1101111;
DRAM[827] = 8'b1101111;
DRAM[828] = 8'b1101111;
DRAM[829] = 8'b1101111;
DRAM[830] = 8'b1101111;
DRAM[831] = 8'b1101111;
DRAM[832] = 8'b1101111;
DRAM[833] = 8'b1101111;
DRAM[834] = 8'b1101111;
DRAM[835] = 8'b1101111;
DRAM[836] = 8'b1101111;
DRAM[837] = 8'b1101110;
DRAM[838] = 8'b1101110;
DRAM[839] = 8'b1101110;
DRAM[840] = 8'b1101110;
DRAM[841] = 8'b1101110;
DRAM[842] = 8'b1101111;
DRAM[843] = 8'b1101111;
DRAM[844] = 8'b1101110;
DRAM[845] = 8'b1101101;
DRAM[846] = 8'b1101100;
DRAM[847] = 8'b1101100;
DRAM[848] = 8'b1101101;
DRAM[849] = 8'b1101101;
DRAM[850] = 8'b1101100;
DRAM[851] = 8'b1101011;
DRAM[852] = 8'b1101011;
DRAM[853] = 8'b1101011;
DRAM[854] = 8'b1101011;
DRAM[855] = 8'b1101011;
DRAM[856] = 8'b1101100;
DRAM[857] = 8'b1101100;
DRAM[858] = 8'b1101100;
DRAM[859] = 8'b1101100;
DRAM[860] = 8'b1101100;
DRAM[861] = 8'b1101100;
DRAM[862] = 8'b1101100;
DRAM[863] = 8'b1101100;
DRAM[864] = 8'b1101011;
DRAM[865] = 8'b1101011;
DRAM[866] = 8'b1101011;
DRAM[867] = 8'b1101011;
DRAM[868] = 8'b1101011;
DRAM[869] = 8'b1101100;
DRAM[870] = 8'b1101101;
DRAM[871] = 8'b1101110;
DRAM[872] = 8'b1101101;
DRAM[873] = 8'b1101100;
DRAM[874] = 8'b1101100;
DRAM[875] = 8'b1101100;
DRAM[876] = 8'b1101011;
DRAM[877] = 8'b1101011;
DRAM[878] = 8'b1101011;
DRAM[879] = 8'b1101011;
DRAM[880] = 8'b1101011;
DRAM[881] = 8'b1101011;
DRAM[882] = 8'b1101011;
DRAM[883] = 8'b1101011;
DRAM[884] = 8'b1101011;
DRAM[885] = 8'b1101011;
DRAM[886] = 8'b1101011;
DRAM[887] = 8'b1101011;
DRAM[888] = 8'b1101010;
DRAM[889] = 8'b1101010;
DRAM[890] = 8'b1101010;
DRAM[891] = 8'b1101010;
DRAM[892] = 8'b1101010;
DRAM[893] = 8'b1101010;
DRAM[894] = 8'b1101010;
DRAM[895] = 8'b1101010;
DRAM[896] = 8'b1101010;
DRAM[897] = 8'b1101010;
DRAM[898] = 8'b1101010;
DRAM[899] = 8'b1101011;
DRAM[900] = 8'b1101011;
DRAM[901] = 8'b1101011;
DRAM[902] = 8'b1101011;
DRAM[903] = 8'b1101011;
DRAM[904] = 8'b1101001;
DRAM[905] = 8'b1101001;
DRAM[906] = 8'b1101010;
DRAM[907] = 8'b1101011;
DRAM[908] = 8'b1101100;
DRAM[909] = 8'b1101100;
DRAM[910] = 8'b1101011;
DRAM[911] = 8'b1101011;
DRAM[912] = 8'b1101000;
DRAM[913] = 8'b1101000;
DRAM[914] = 8'b1101001;
DRAM[915] = 8'b1101001;
DRAM[916] = 8'b1101001;
DRAM[917] = 8'b1101001;
DRAM[918] = 8'b1101000;
DRAM[919] = 8'b1101000;
DRAM[920] = 8'b1100111;
DRAM[921] = 8'b1100111;
DRAM[922] = 8'b1100111;
DRAM[923] = 8'b1100111;
DRAM[924] = 8'b1100111;
DRAM[925] = 8'b1100111;
DRAM[926] = 8'b1100111;
DRAM[927] = 8'b1100111;
DRAM[928] = 8'b1101000;
DRAM[929] = 8'b1101000;
DRAM[930] = 8'b1101000;
DRAM[931] = 8'b1101000;
DRAM[932] = 8'b1100111;
DRAM[933] = 8'b1100110;
DRAM[934] = 8'b1100100;
DRAM[935] = 8'b1100100;
DRAM[936] = 8'b1100100;
DRAM[937] = 8'b1100100;
DRAM[938] = 8'b1100011;
DRAM[939] = 8'b1100010;
DRAM[940] = 8'b1100010;
DRAM[941] = 8'b1100010;
DRAM[942] = 8'b1100010;
DRAM[943] = 8'b1100010;
DRAM[944] = 8'b1100001;
DRAM[945] = 8'b1100000;
DRAM[946] = 8'b1100000;
DRAM[947] = 8'b1100000;
DRAM[948] = 8'b1011111;
DRAM[949] = 8'b1011111;
DRAM[950] = 8'b1011111;
DRAM[951] = 8'b1011111;
DRAM[952] = 8'b1011101;
DRAM[953] = 8'b1011101;
DRAM[954] = 8'b1011101;
DRAM[955] = 8'b1011100;
DRAM[956] = 8'b1011011;
DRAM[957] = 8'b1011010;
DRAM[958] = 8'b1011010;
DRAM[959] = 8'b1011001;
DRAM[960] = 8'b1010111;
DRAM[961] = 8'b1010111;
DRAM[962] = 8'b1010111;
DRAM[963] = 8'b1010111;
DRAM[964] = 8'b1010110;
DRAM[965] = 8'b1010110;
DRAM[966] = 8'b1010110;
DRAM[967] = 8'b1010110;
DRAM[968] = 8'b1010101;
DRAM[969] = 8'b1010100;
DRAM[970] = 8'b1010100;
DRAM[971] = 8'b1010100;
DRAM[972] = 8'b1010011;
DRAM[973] = 8'b1010011;
DRAM[974] = 8'b1010011;
DRAM[975] = 8'b1010011;
DRAM[976] = 8'b1010001;
DRAM[977] = 8'b1010001;
DRAM[978] = 8'b1010000;
DRAM[979] = 8'b1010000;
DRAM[980] = 8'b1010000;
DRAM[981] = 8'b1001111;
DRAM[982] = 8'b1001111;
DRAM[983] = 8'b1001111;
DRAM[984] = 8'b1010001;
DRAM[985] = 8'b1010001;
DRAM[986] = 8'b1010000;
DRAM[987] = 8'b1001111;
DRAM[988] = 8'b1001110;
DRAM[989] = 8'b1001100;
DRAM[990] = 8'b1001010;
DRAM[991] = 8'b1001001;
DRAM[992] = 8'b1001001;
DRAM[993] = 8'b1001000;
DRAM[994] = 8'b1001000;
DRAM[995] = 8'b1001000;
DRAM[996] = 8'b1000111;
DRAM[997] = 8'b1000111;
DRAM[998] = 8'b1000111;
DRAM[999] = 8'b1000111;
DRAM[1000] = 8'b1000111;
DRAM[1001] = 8'b1000110;
DRAM[1002] = 8'b1000110;
DRAM[1003] = 8'b1000110;
DRAM[1004] = 8'b1000101;
DRAM[1005] = 8'b1000101;
DRAM[1006] = 8'b1000101;
DRAM[1007] = 8'b1000100;
DRAM[1008] = 8'b1000011;
DRAM[1009] = 8'b1000011;
DRAM[1010] = 8'b1000010;
DRAM[1011] = 8'b1000010;
DRAM[1012] = 8'b1000010;
DRAM[1013] = 8'b1000001;
DRAM[1014] = 8'b1000001;
DRAM[1015] = 8'b1000001;
DRAM[1016] = 8'b111111;
DRAM[1017] = 8'b111111;
DRAM[1018] = 8'b111110;
DRAM[1019] = 8'b111110;
DRAM[1020] = 8'b111101;
DRAM[1021] = 8'b111101;
DRAM[1022] = 8'b111101;
DRAM[1023] = 8'b111101;
DRAM[1024] = 8'b1011010;
DRAM[1025] = 8'b1011011;
DRAM[1026] = 8'b1011011;
DRAM[1027] = 8'b1011100;
DRAM[1028] = 8'b1011101;
DRAM[1029] = 8'b1011110;
DRAM[1030] = 8'b1011110;
DRAM[1031] = 8'b1011110;
DRAM[1032] = 8'b1011110;
DRAM[1033] = 8'b1011101;
DRAM[1034] = 8'b1011101;
DRAM[1035] = 8'b1011111;
DRAM[1036] = 8'b1100010;
DRAM[1037] = 8'b1100100;
DRAM[1038] = 8'b1100011;
DRAM[1039] = 8'b1100010;
DRAM[1040] = 8'b1100110;
DRAM[1041] = 8'b1100101;
DRAM[1042] = 8'b1100100;
DRAM[1043] = 8'b1100100;
DRAM[1044] = 8'b1100100;
DRAM[1045] = 8'b1100110;
DRAM[1046] = 8'b1100111;
DRAM[1047] = 8'b1101000;
DRAM[1048] = 8'b1100110;
DRAM[1049] = 8'b1100110;
DRAM[1050] = 8'b1100110;
DRAM[1051] = 8'b1100111;
DRAM[1052] = 8'b1100111;
DRAM[1053] = 8'b1100111;
DRAM[1054] = 8'b1101000;
DRAM[1055] = 8'b1101000;
DRAM[1056] = 8'b1100111;
DRAM[1057] = 8'b1100111;
DRAM[1058] = 8'b1101000;
DRAM[1059] = 8'b1101001;
DRAM[1060] = 8'b1101010;
DRAM[1061] = 8'b1101011;
DRAM[1062] = 8'b1101011;
DRAM[1063] = 8'b1101100;
DRAM[1064] = 8'b1101100;
DRAM[1065] = 8'b1101100;
DRAM[1066] = 8'b1101101;
DRAM[1067] = 8'b1101101;
DRAM[1068] = 8'b1101110;
DRAM[1069] = 8'b1101110;
DRAM[1070] = 8'b1101111;
DRAM[1071] = 8'b1101111;
DRAM[1072] = 8'b1101110;
DRAM[1073] = 8'b1101110;
DRAM[1074] = 8'b1101110;
DRAM[1075] = 8'b1101110;
DRAM[1076] = 8'b1101110;
DRAM[1077] = 8'b1101110;
DRAM[1078] = 8'b1101110;
DRAM[1079] = 8'b1101110;
DRAM[1080] = 8'b1101111;
DRAM[1081] = 8'b1101111;
DRAM[1082] = 8'b1101111;
DRAM[1083] = 8'b1101111;
DRAM[1084] = 8'b1101111;
DRAM[1085] = 8'b1101111;
DRAM[1086] = 8'b1101111;
DRAM[1087] = 8'b1101111;
DRAM[1088] = 8'b1101111;
DRAM[1089] = 8'b1101111;
DRAM[1090] = 8'b1101111;
DRAM[1091] = 8'b1101111;
DRAM[1092] = 8'b1101111;
DRAM[1093] = 8'b1110000;
DRAM[1094] = 8'b1110000;
DRAM[1095] = 8'b1110000;
DRAM[1096] = 8'b1101111;
DRAM[1097] = 8'b1101111;
DRAM[1098] = 8'b1101111;
DRAM[1099] = 8'b1101111;
DRAM[1100] = 8'b1101111;
DRAM[1101] = 8'b1101110;
DRAM[1102] = 8'b1101101;
DRAM[1103] = 8'b1101101;
DRAM[1104] = 8'b1101110;
DRAM[1105] = 8'b1101110;
DRAM[1106] = 8'b1101101;
DRAM[1107] = 8'b1101100;
DRAM[1108] = 8'b1101011;
DRAM[1109] = 8'b1101011;
DRAM[1110] = 8'b1101100;
DRAM[1111] = 8'b1101100;
DRAM[1112] = 8'b1101100;
DRAM[1113] = 8'b1101100;
DRAM[1114] = 8'b1101100;
DRAM[1115] = 8'b1101100;
DRAM[1116] = 8'b1101100;
DRAM[1117] = 8'b1101100;
DRAM[1118] = 8'b1101100;
DRAM[1119] = 8'b1101100;
DRAM[1120] = 8'b1101100;
DRAM[1121] = 8'b1101100;
DRAM[1122] = 8'b1101011;
DRAM[1123] = 8'b1101011;
DRAM[1124] = 8'b1101011;
DRAM[1125] = 8'b1101100;
DRAM[1126] = 8'b1101101;
DRAM[1127] = 8'b1101110;
DRAM[1128] = 8'b1101101;
DRAM[1129] = 8'b1101101;
DRAM[1130] = 8'b1101101;
DRAM[1131] = 8'b1101101;
DRAM[1132] = 8'b1101100;
DRAM[1133] = 8'b1101100;
DRAM[1134] = 8'b1101100;
DRAM[1135] = 8'b1101011;
DRAM[1136] = 8'b1101011;
DRAM[1137] = 8'b1101011;
DRAM[1138] = 8'b1101011;
DRAM[1139] = 8'b1101011;
DRAM[1140] = 8'b1101011;
DRAM[1141] = 8'b1101011;
DRAM[1142] = 8'b1101011;
DRAM[1143] = 8'b1101011;
DRAM[1144] = 8'b1101010;
DRAM[1145] = 8'b1101010;
DRAM[1146] = 8'b1101010;
DRAM[1147] = 8'b1101010;
DRAM[1148] = 8'b1101010;
DRAM[1149] = 8'b1101010;
DRAM[1150] = 8'b1101010;
DRAM[1151] = 8'b1101010;
DRAM[1152] = 8'b1101100;
DRAM[1153] = 8'b1101100;
DRAM[1154] = 8'b1101100;
DRAM[1155] = 8'b1101011;
DRAM[1156] = 8'b1101011;
DRAM[1157] = 8'b1101011;
DRAM[1158] = 8'b1101011;
DRAM[1159] = 8'b1101011;
DRAM[1160] = 8'b1101010;
DRAM[1161] = 8'b1101010;
DRAM[1162] = 8'b1101011;
DRAM[1163] = 8'b1101100;
DRAM[1164] = 8'b1101100;
DRAM[1165] = 8'b1101100;
DRAM[1166] = 8'b1101100;
DRAM[1167] = 8'b1101100;
DRAM[1168] = 8'b1101010;
DRAM[1169] = 8'b1101011;
DRAM[1170] = 8'b1101011;
DRAM[1171] = 8'b1101100;
DRAM[1172] = 8'b1101100;
DRAM[1173] = 8'b1101011;
DRAM[1174] = 8'b1101011;
DRAM[1175] = 8'b1101010;
DRAM[1176] = 8'b1101001;
DRAM[1177] = 8'b1101001;
DRAM[1178] = 8'b1101001;
DRAM[1179] = 8'b1101001;
DRAM[1180] = 8'b1101001;
DRAM[1181] = 8'b1101001;
DRAM[1182] = 8'b1101001;
DRAM[1183] = 8'b1101001;
DRAM[1184] = 8'b1101001;
DRAM[1185] = 8'b1101001;
DRAM[1186] = 8'b1101001;
DRAM[1187] = 8'b1101001;
DRAM[1188] = 8'b1101000;
DRAM[1189] = 8'b1100111;
DRAM[1190] = 8'b1100101;
DRAM[1191] = 8'b1100101;
DRAM[1192] = 8'b1100100;
DRAM[1193] = 8'b1100100;
DRAM[1194] = 8'b1100100;
DRAM[1195] = 8'b1100100;
DRAM[1196] = 8'b1100100;
DRAM[1197] = 8'b1100011;
DRAM[1198] = 8'b1100010;
DRAM[1199] = 8'b1100010;
DRAM[1200] = 8'b1100001;
DRAM[1201] = 8'b1100001;
DRAM[1202] = 8'b1100001;
DRAM[1203] = 8'b1100001;
DRAM[1204] = 8'b1100000;
DRAM[1205] = 8'b1100000;
DRAM[1206] = 8'b1100000;
DRAM[1207] = 8'b1011111;
DRAM[1208] = 8'b1011111;
DRAM[1209] = 8'b1011110;
DRAM[1210] = 8'b1011110;
DRAM[1211] = 8'b1011101;
DRAM[1212] = 8'b1011100;
DRAM[1213] = 8'b1011011;
DRAM[1214] = 8'b1011011;
DRAM[1215] = 8'b1011011;
DRAM[1216] = 8'b1011001;
DRAM[1217] = 8'b1011001;
DRAM[1218] = 8'b1011000;
DRAM[1219] = 8'b1011000;
DRAM[1220] = 8'b1010111;
DRAM[1221] = 8'b1010111;
DRAM[1222] = 8'b1010110;
DRAM[1223] = 8'b1010110;
DRAM[1224] = 8'b1010101;
DRAM[1225] = 8'b1010101;
DRAM[1226] = 8'b1010101;
DRAM[1227] = 8'b1010101;
DRAM[1228] = 8'b1010100;
DRAM[1229] = 8'b1010100;
DRAM[1230] = 8'b1010100;
DRAM[1231] = 8'b1010011;
DRAM[1232] = 8'b1010001;
DRAM[1233] = 8'b1010001;
DRAM[1234] = 8'b1010001;
DRAM[1235] = 8'b1010000;
DRAM[1236] = 8'b1010000;
DRAM[1237] = 8'b1010000;
DRAM[1238] = 8'b1001111;
DRAM[1239] = 8'b1001111;
DRAM[1240] = 8'b1010001;
DRAM[1241] = 8'b1010001;
DRAM[1242] = 8'b1010001;
DRAM[1243] = 8'b1010000;
DRAM[1244] = 8'b1001111;
DRAM[1245] = 8'b1001101;
DRAM[1246] = 8'b1001011;
DRAM[1247] = 8'b1001010;
DRAM[1248] = 8'b1001001;
DRAM[1249] = 8'b1001001;
DRAM[1250] = 8'b1001001;
DRAM[1251] = 8'b1001001;
DRAM[1252] = 8'b1001000;
DRAM[1253] = 8'b1001000;
DRAM[1254] = 8'b1001000;
DRAM[1255] = 8'b1000111;
DRAM[1256] = 8'b1000110;
DRAM[1257] = 8'b1000101;
DRAM[1258] = 8'b1000101;
DRAM[1259] = 8'b1000101;
DRAM[1260] = 8'b1000100;
DRAM[1261] = 8'b1000100;
DRAM[1262] = 8'b1000100;
DRAM[1263] = 8'b1000011;
DRAM[1264] = 8'b1000011;
DRAM[1265] = 8'b1000011;
DRAM[1266] = 8'b1000011;
DRAM[1267] = 8'b1000010;
DRAM[1268] = 8'b1000010;
DRAM[1269] = 8'b1000010;
DRAM[1270] = 8'b1000001;
DRAM[1271] = 8'b1000001;
DRAM[1272] = 8'b111111;
DRAM[1273] = 8'b111111;
DRAM[1274] = 8'b111111;
DRAM[1275] = 8'b111110;
DRAM[1276] = 8'b111110;
DRAM[1277] = 8'b111101;
DRAM[1278] = 8'b111101;
DRAM[1279] = 8'b111101;
DRAM[1280] = 8'b1011011;
DRAM[1281] = 8'b1011011;
DRAM[1282] = 8'b1011100;
DRAM[1283] = 8'b1011101;
DRAM[1284] = 8'b1011110;
DRAM[1285] = 8'b1011110;
DRAM[1286] = 8'b1011111;
DRAM[1287] = 8'b1011111;
DRAM[1288] = 8'b1011111;
DRAM[1289] = 8'b1011110;
DRAM[1290] = 8'b1011110;
DRAM[1291] = 8'b1100000;
DRAM[1292] = 8'b1100011;
DRAM[1293] = 8'b1100100;
DRAM[1294] = 8'b1100100;
DRAM[1295] = 8'b1100011;
DRAM[1296] = 8'b1100110;
DRAM[1297] = 8'b1100110;
DRAM[1298] = 8'b1100110;
DRAM[1299] = 8'b1100110;
DRAM[1300] = 8'b1100110;
DRAM[1301] = 8'b1100111;
DRAM[1302] = 8'b1101000;
DRAM[1303] = 8'b1101001;
DRAM[1304] = 8'b1100111;
DRAM[1305] = 8'b1100111;
DRAM[1306] = 8'b1100111;
DRAM[1307] = 8'b1101000;
DRAM[1308] = 8'b1101000;
DRAM[1309] = 8'b1101000;
DRAM[1310] = 8'b1101001;
DRAM[1311] = 8'b1101001;
DRAM[1312] = 8'b1100111;
DRAM[1313] = 8'b1101000;
DRAM[1314] = 8'b1101001;
DRAM[1315] = 8'b1101010;
DRAM[1316] = 8'b1101011;
DRAM[1317] = 8'b1101100;
DRAM[1318] = 8'b1101101;
DRAM[1319] = 8'b1101101;
DRAM[1320] = 8'b1101100;
DRAM[1321] = 8'b1101101;
DRAM[1322] = 8'b1101101;
DRAM[1323] = 8'b1101110;
DRAM[1324] = 8'b1101111;
DRAM[1325] = 8'b1101111;
DRAM[1326] = 8'b1110000;
DRAM[1327] = 8'b1110000;
DRAM[1328] = 8'b1101111;
DRAM[1329] = 8'b1101111;
DRAM[1330] = 8'b1101111;
DRAM[1331] = 8'b1101111;
DRAM[1332] = 8'b1101111;
DRAM[1333] = 8'b1101111;
DRAM[1334] = 8'b1101111;
DRAM[1335] = 8'b1101111;
DRAM[1336] = 8'b1110000;
DRAM[1337] = 8'b1110000;
DRAM[1338] = 8'b1110000;
DRAM[1339] = 8'b1110000;
DRAM[1340] = 8'b1110000;
DRAM[1341] = 8'b1110000;
DRAM[1342] = 8'b1110000;
DRAM[1343] = 8'b1110000;
DRAM[1344] = 8'b1101111;
DRAM[1345] = 8'b1101111;
DRAM[1346] = 8'b1110000;
DRAM[1347] = 8'b1110000;
DRAM[1348] = 8'b1110000;
DRAM[1349] = 8'b1110001;
DRAM[1350] = 8'b1110001;
DRAM[1351] = 8'b1110001;
DRAM[1352] = 8'b1101111;
DRAM[1353] = 8'b1110000;
DRAM[1354] = 8'b1110000;
DRAM[1355] = 8'b1110000;
DRAM[1356] = 8'b1110000;
DRAM[1357] = 8'b1101111;
DRAM[1358] = 8'b1101110;
DRAM[1359] = 8'b1101101;
DRAM[1360] = 8'b1101111;
DRAM[1361] = 8'b1101110;
DRAM[1362] = 8'b1101101;
DRAM[1363] = 8'b1101101;
DRAM[1364] = 8'b1101100;
DRAM[1365] = 8'b1101100;
DRAM[1366] = 8'b1101101;
DRAM[1367] = 8'b1101101;
DRAM[1368] = 8'b1101101;
DRAM[1369] = 8'b1101101;
DRAM[1370] = 8'b1101101;
DRAM[1371] = 8'b1101101;
DRAM[1372] = 8'b1101101;
DRAM[1373] = 8'b1101101;
DRAM[1374] = 8'b1101101;
DRAM[1375] = 8'b1101101;
DRAM[1376] = 8'b1101101;
DRAM[1377] = 8'b1101101;
DRAM[1378] = 8'b1101100;
DRAM[1379] = 8'b1101100;
DRAM[1380] = 8'b1101101;
DRAM[1381] = 8'b1101101;
DRAM[1382] = 8'b1101110;
DRAM[1383] = 8'b1101111;
DRAM[1384] = 8'b1101110;
DRAM[1385] = 8'b1101110;
DRAM[1386] = 8'b1101110;
DRAM[1387] = 8'b1101101;
DRAM[1388] = 8'b1101101;
DRAM[1389] = 8'b1101101;
DRAM[1390] = 8'b1101100;
DRAM[1391] = 8'b1101100;
DRAM[1392] = 8'b1101100;
DRAM[1393] = 8'b1101100;
DRAM[1394] = 8'b1101100;
DRAM[1395] = 8'b1101100;
DRAM[1396] = 8'b1101100;
DRAM[1397] = 8'b1101100;
DRAM[1398] = 8'b1101100;
DRAM[1399] = 8'b1101100;
DRAM[1400] = 8'b1101011;
DRAM[1401] = 8'b1101011;
DRAM[1402] = 8'b1101011;
DRAM[1403] = 8'b1101011;
DRAM[1404] = 8'b1101011;
DRAM[1405] = 8'b1101011;
DRAM[1406] = 8'b1101011;
DRAM[1407] = 8'b1101011;
DRAM[1408] = 8'b1101101;
DRAM[1409] = 8'b1101101;
DRAM[1410] = 8'b1101101;
DRAM[1411] = 8'b1101100;
DRAM[1412] = 8'b1101100;
DRAM[1413] = 8'b1101100;
DRAM[1414] = 8'b1101011;
DRAM[1415] = 8'b1101011;
DRAM[1416] = 8'b1101010;
DRAM[1417] = 8'b1101011;
DRAM[1418] = 8'b1101100;
DRAM[1419] = 8'b1101101;
DRAM[1420] = 8'b1101101;
DRAM[1421] = 8'b1101101;
DRAM[1422] = 8'b1101101;
DRAM[1423] = 8'b1101100;
DRAM[1424] = 8'b1101101;
DRAM[1425] = 8'b1101101;
DRAM[1426] = 8'b1101110;
DRAM[1427] = 8'b1101110;
DRAM[1428] = 8'b1101110;
DRAM[1429] = 8'b1101110;
DRAM[1430] = 8'b1101101;
DRAM[1431] = 8'b1101101;
DRAM[1432] = 8'b1101100;
DRAM[1433] = 8'b1101100;
DRAM[1434] = 8'b1101100;
DRAM[1435] = 8'b1101100;
DRAM[1436] = 8'b1101100;
DRAM[1437] = 8'b1101100;
DRAM[1438] = 8'b1101100;
DRAM[1439] = 8'b1101100;
DRAM[1440] = 8'b1101001;
DRAM[1441] = 8'b1101010;
DRAM[1442] = 8'b1101010;
DRAM[1443] = 8'b1101001;
DRAM[1444] = 8'b1101001;
DRAM[1445] = 8'b1100111;
DRAM[1446] = 8'b1100110;
DRAM[1447] = 8'b1100101;
DRAM[1448] = 8'b1100100;
DRAM[1449] = 8'b1100101;
DRAM[1450] = 8'b1100101;
DRAM[1451] = 8'b1100101;
DRAM[1452] = 8'b1100101;
DRAM[1453] = 8'b1100100;
DRAM[1454] = 8'b1100011;
DRAM[1455] = 8'b1100010;
DRAM[1456] = 8'b1100010;
DRAM[1457] = 8'b1100010;
DRAM[1458] = 8'b1100010;
DRAM[1459] = 8'b1100001;
DRAM[1460] = 8'b1100001;
DRAM[1461] = 8'b1100001;
DRAM[1462] = 8'b1100000;
DRAM[1463] = 8'b1100000;
DRAM[1464] = 8'b1100000;
DRAM[1465] = 8'b1100000;
DRAM[1466] = 8'b1011111;
DRAM[1467] = 8'b1011110;
DRAM[1468] = 8'b1011101;
DRAM[1469] = 8'b1011101;
DRAM[1470] = 8'b1011100;
DRAM[1471] = 8'b1011100;
DRAM[1472] = 8'b1011010;
DRAM[1473] = 8'b1011010;
DRAM[1474] = 8'b1011001;
DRAM[1475] = 8'b1011001;
DRAM[1476] = 8'b1011000;
DRAM[1477] = 8'b1010111;
DRAM[1478] = 8'b1010111;
DRAM[1479] = 8'b1010110;
DRAM[1480] = 8'b1010110;
DRAM[1481] = 8'b1010110;
DRAM[1482] = 8'b1010110;
DRAM[1483] = 8'b1010101;
DRAM[1484] = 8'b1010101;
DRAM[1485] = 8'b1010101;
DRAM[1486] = 8'b1010100;
DRAM[1487] = 8'b1010100;
DRAM[1488] = 8'b1010010;
DRAM[1489] = 8'b1010001;
DRAM[1490] = 8'b1010001;
DRAM[1491] = 8'b1010001;
DRAM[1492] = 8'b1010000;
DRAM[1493] = 8'b1010000;
DRAM[1494] = 8'b1010000;
DRAM[1495] = 8'b1010000;
DRAM[1496] = 8'b1010001;
DRAM[1497] = 8'b1010001;
DRAM[1498] = 8'b1010001;
DRAM[1499] = 8'b1010000;
DRAM[1500] = 8'b1001111;
DRAM[1501] = 8'b1001101;
DRAM[1502] = 8'b1001100;
DRAM[1503] = 8'b1001011;
DRAM[1504] = 8'b1001010;
DRAM[1505] = 8'b1001010;
DRAM[1506] = 8'b1001010;
DRAM[1507] = 8'b1001001;
DRAM[1508] = 8'b1001001;
DRAM[1509] = 8'b1001001;
DRAM[1510] = 8'b1001000;
DRAM[1511] = 8'b1001000;
DRAM[1512] = 8'b1000101;
DRAM[1513] = 8'b1000101;
DRAM[1514] = 8'b1000101;
DRAM[1515] = 8'b1000101;
DRAM[1516] = 8'b1000100;
DRAM[1517] = 8'b1000100;
DRAM[1518] = 8'b1000011;
DRAM[1519] = 8'b1000011;
DRAM[1520] = 8'b1000100;
DRAM[1521] = 8'b1000011;
DRAM[1522] = 8'b1000011;
DRAM[1523] = 8'b1000011;
DRAM[1524] = 8'b1000010;
DRAM[1525] = 8'b1000010;
DRAM[1526] = 8'b1000010;
DRAM[1527] = 8'b1000010;
DRAM[1528] = 8'b1000000;
DRAM[1529] = 8'b1000000;
DRAM[1530] = 8'b1000000;
DRAM[1531] = 8'b111111;
DRAM[1532] = 8'b111111;
DRAM[1533] = 8'b111111;
DRAM[1534] = 8'b111110;
DRAM[1535] = 8'b111110;
DRAM[1536] = 8'b1011100;
DRAM[1537] = 8'b1011100;
DRAM[1538] = 8'b1011101;
DRAM[1539] = 8'b1011101;
DRAM[1540] = 8'b1011110;
DRAM[1541] = 8'b1011111;
DRAM[1542] = 8'b1100000;
DRAM[1543] = 8'b1100000;
DRAM[1544] = 8'b1100000;
DRAM[1545] = 8'b1011111;
DRAM[1546] = 8'b1011111;
DRAM[1547] = 8'b1100000;
DRAM[1548] = 8'b1100011;
DRAM[1549] = 8'b1100101;
DRAM[1550] = 8'b1100101;
DRAM[1551] = 8'b1100100;
DRAM[1552] = 8'b1100110;
DRAM[1553] = 8'b1100110;
DRAM[1554] = 8'b1100111;
DRAM[1555] = 8'b1101000;
DRAM[1556] = 8'b1101001;
DRAM[1557] = 8'b1101001;
DRAM[1558] = 8'b1101000;
DRAM[1559] = 8'b1101000;
DRAM[1560] = 8'b1100110;
DRAM[1561] = 8'b1100110;
DRAM[1562] = 8'b1100111;
DRAM[1563] = 8'b1100111;
DRAM[1564] = 8'b1100111;
DRAM[1565] = 8'b1101000;
DRAM[1566] = 8'b1101000;
DRAM[1567] = 8'b1101000;
DRAM[1568] = 8'b1100111;
DRAM[1569] = 8'b1101000;
DRAM[1570] = 8'b1101001;
DRAM[1571] = 8'b1101010;
DRAM[1572] = 8'b1101011;
DRAM[1573] = 8'b1101101;
DRAM[1574] = 8'b1101110;
DRAM[1575] = 8'b1101110;
DRAM[1576] = 8'b1101100;
DRAM[1577] = 8'b1101101;
DRAM[1578] = 8'b1101101;
DRAM[1579] = 8'b1101110;
DRAM[1580] = 8'b1101111;
DRAM[1581] = 8'b1110000;
DRAM[1582] = 8'b1110001;
DRAM[1583] = 8'b1110001;
DRAM[1584] = 8'b1110000;
DRAM[1585] = 8'b1110000;
DRAM[1586] = 8'b1110000;
DRAM[1587] = 8'b1110000;
DRAM[1588] = 8'b1110000;
DRAM[1589] = 8'b1110000;
DRAM[1590] = 8'b1110000;
DRAM[1591] = 8'b1110000;
DRAM[1592] = 8'b1110001;
DRAM[1593] = 8'b1110001;
DRAM[1594] = 8'b1110001;
DRAM[1595] = 8'b1110001;
DRAM[1596] = 8'b1110001;
DRAM[1597] = 8'b1110001;
DRAM[1598] = 8'b1110001;
DRAM[1599] = 8'b1110001;
DRAM[1600] = 8'b1110000;
DRAM[1601] = 8'b1110000;
DRAM[1602] = 8'b1110000;
DRAM[1603] = 8'b1110001;
DRAM[1604] = 8'b1110001;
DRAM[1605] = 8'b1110001;
DRAM[1606] = 8'b1110010;
DRAM[1607] = 8'b1110010;
DRAM[1608] = 8'b1110000;
DRAM[1609] = 8'b1110000;
DRAM[1610] = 8'b1110001;
DRAM[1611] = 8'b1110001;
DRAM[1612] = 8'b1110000;
DRAM[1613] = 8'b1101111;
DRAM[1614] = 8'b1101111;
DRAM[1615] = 8'b1101110;
DRAM[1616] = 8'b1110000;
DRAM[1617] = 8'b1101111;
DRAM[1618] = 8'b1101110;
DRAM[1619] = 8'b1101101;
DRAM[1620] = 8'b1101101;
DRAM[1621] = 8'b1101101;
DRAM[1622] = 8'b1101101;
DRAM[1623] = 8'b1101110;
DRAM[1624] = 8'b1101110;
DRAM[1625] = 8'b1101110;
DRAM[1626] = 8'b1101110;
DRAM[1627] = 8'b1101110;
DRAM[1628] = 8'b1101110;
DRAM[1629] = 8'b1101110;
DRAM[1630] = 8'b1101110;
DRAM[1631] = 8'b1101110;
DRAM[1632] = 8'b1101110;
DRAM[1633] = 8'b1101110;
DRAM[1634] = 8'b1101101;
DRAM[1635] = 8'b1101101;
DRAM[1636] = 8'b1101110;
DRAM[1637] = 8'b1101111;
DRAM[1638] = 8'b1110000;
DRAM[1639] = 8'b1110000;
DRAM[1640] = 8'b1101111;
DRAM[1641] = 8'b1101111;
DRAM[1642] = 8'b1101110;
DRAM[1643] = 8'b1101110;
DRAM[1644] = 8'b1101110;
DRAM[1645] = 8'b1101101;
DRAM[1646] = 8'b1101101;
DRAM[1647] = 8'b1101101;
DRAM[1648] = 8'b1101101;
DRAM[1649] = 8'b1101101;
DRAM[1650] = 8'b1101101;
DRAM[1651] = 8'b1101101;
DRAM[1652] = 8'b1101101;
DRAM[1653] = 8'b1101101;
DRAM[1654] = 8'b1101101;
DRAM[1655] = 8'b1101101;
DRAM[1656] = 8'b1101100;
DRAM[1657] = 8'b1101100;
DRAM[1658] = 8'b1101100;
DRAM[1659] = 8'b1101100;
DRAM[1660] = 8'b1101100;
DRAM[1661] = 8'b1101100;
DRAM[1662] = 8'b1101100;
DRAM[1663] = 8'b1101100;
DRAM[1664] = 8'b1101110;
DRAM[1665] = 8'b1101110;
DRAM[1666] = 8'b1101101;
DRAM[1667] = 8'b1101101;
DRAM[1668] = 8'b1101101;
DRAM[1669] = 8'b1101100;
DRAM[1670] = 8'b1101100;
DRAM[1671] = 8'b1101100;
DRAM[1672] = 8'b1101011;
DRAM[1673] = 8'b1101100;
DRAM[1674] = 8'b1101100;
DRAM[1675] = 8'b1101101;
DRAM[1676] = 8'b1101110;
DRAM[1677] = 8'b1101110;
DRAM[1678] = 8'b1101101;
DRAM[1679] = 8'b1101101;
DRAM[1680] = 8'b1101110;
DRAM[1681] = 8'b1101110;
DRAM[1682] = 8'b1101111;
DRAM[1683] = 8'b1101111;
DRAM[1684] = 8'b1101111;
DRAM[1685] = 8'b1101111;
DRAM[1686] = 8'b1101110;
DRAM[1687] = 8'b1101110;
DRAM[1688] = 8'b1101100;
DRAM[1689] = 8'b1101100;
DRAM[1690] = 8'b1101100;
DRAM[1691] = 8'b1101100;
DRAM[1692] = 8'b1101100;
DRAM[1693] = 8'b1101100;
DRAM[1694] = 8'b1101100;
DRAM[1695] = 8'b1101100;
DRAM[1696] = 8'b1101010;
DRAM[1697] = 8'b1101010;
DRAM[1698] = 8'b1101010;
DRAM[1699] = 8'b1101010;
DRAM[1700] = 8'b1101001;
DRAM[1701] = 8'b1101000;
DRAM[1702] = 8'b1100111;
DRAM[1703] = 8'b1100110;
DRAM[1704] = 8'b1100100;
DRAM[1705] = 8'b1100101;
DRAM[1706] = 8'b1100110;
DRAM[1707] = 8'b1100110;
DRAM[1708] = 8'b1100110;
DRAM[1709] = 8'b1100101;
DRAM[1710] = 8'b1100011;
DRAM[1711] = 8'b1100010;
DRAM[1712] = 8'b1100011;
DRAM[1713] = 8'b1100011;
DRAM[1714] = 8'b1100010;
DRAM[1715] = 8'b1100010;
DRAM[1716] = 8'b1100010;
DRAM[1717] = 8'b1100001;
DRAM[1718] = 8'b1100001;
DRAM[1719] = 8'b1100001;
DRAM[1720] = 8'b1100001;
DRAM[1721] = 8'b1100000;
DRAM[1722] = 8'b1100000;
DRAM[1723] = 8'b1011111;
DRAM[1724] = 8'b1011110;
DRAM[1725] = 8'b1011101;
DRAM[1726] = 8'b1011101;
DRAM[1727] = 8'b1011101;
DRAM[1728] = 8'b1011011;
DRAM[1729] = 8'b1011011;
DRAM[1730] = 8'b1011010;
DRAM[1731] = 8'b1011001;
DRAM[1732] = 8'b1011000;
DRAM[1733] = 8'b1010111;
DRAM[1734] = 8'b1010111;
DRAM[1735] = 8'b1010110;
DRAM[1736] = 8'b1010111;
DRAM[1737] = 8'b1010111;
DRAM[1738] = 8'b1010110;
DRAM[1739] = 8'b1010110;
DRAM[1740] = 8'b1010110;
DRAM[1741] = 8'b1010101;
DRAM[1742] = 8'b1010101;
DRAM[1743] = 8'b1010101;
DRAM[1744] = 8'b1010010;
DRAM[1745] = 8'b1010010;
DRAM[1746] = 8'b1010001;
DRAM[1747] = 8'b1010001;
DRAM[1748] = 8'b1010001;
DRAM[1749] = 8'b1010000;
DRAM[1750] = 8'b1010000;
DRAM[1751] = 8'b1010000;
DRAM[1752] = 8'b1001111;
DRAM[1753] = 8'b1001111;
DRAM[1754] = 8'b1001111;
DRAM[1755] = 8'b1001111;
DRAM[1756] = 8'b1001111;
DRAM[1757] = 8'b1001110;
DRAM[1758] = 8'b1001101;
DRAM[1759] = 8'b1001100;
DRAM[1760] = 8'b1001011;
DRAM[1761] = 8'b1001011;
DRAM[1762] = 8'b1001010;
DRAM[1763] = 8'b1001010;
DRAM[1764] = 8'b1001010;
DRAM[1765] = 8'b1001001;
DRAM[1766] = 8'b1001001;
DRAM[1767] = 8'b1001001;
DRAM[1768] = 8'b1000111;
DRAM[1769] = 8'b1000111;
DRAM[1770] = 8'b1000110;
DRAM[1771] = 8'b1000110;
DRAM[1772] = 8'b1000101;
DRAM[1773] = 8'b1000101;
DRAM[1774] = 8'b1000101;
DRAM[1775] = 8'b1000101;
DRAM[1776] = 8'b1000100;
DRAM[1777] = 8'b1000100;
DRAM[1778] = 8'b1000011;
DRAM[1779] = 8'b1000011;
DRAM[1780] = 8'b1000011;
DRAM[1781] = 8'b1000010;
DRAM[1782] = 8'b1000010;
DRAM[1783] = 8'b1000010;
DRAM[1784] = 8'b1000001;
DRAM[1785] = 8'b1000001;
DRAM[1786] = 8'b1000001;
DRAM[1787] = 8'b1000001;
DRAM[1788] = 8'b1000000;
DRAM[1789] = 8'b1000000;
DRAM[1790] = 8'b111111;
DRAM[1791] = 8'b111111;
DRAM[1792] = 8'b1011100;
DRAM[1793] = 8'b1011100;
DRAM[1794] = 8'b1011101;
DRAM[1795] = 8'b1011110;
DRAM[1796] = 8'b1011111;
DRAM[1797] = 8'b1011111;
DRAM[1798] = 8'b1100000;
DRAM[1799] = 8'b1100000;
DRAM[1800] = 8'b1100000;
DRAM[1801] = 8'b1011111;
DRAM[1802] = 8'b1011111;
DRAM[1803] = 8'b1100001;
DRAM[1804] = 8'b1100100;
DRAM[1805] = 8'b1100101;
DRAM[1806] = 8'b1100101;
DRAM[1807] = 8'b1100100;
DRAM[1808] = 8'b1100101;
DRAM[1809] = 8'b1100111;
DRAM[1810] = 8'b1101000;
DRAM[1811] = 8'b1101010;
DRAM[1812] = 8'b1101010;
DRAM[1813] = 8'b1101001;
DRAM[1814] = 8'b1101000;
DRAM[1815] = 8'b1100111;
DRAM[1816] = 8'b1100101;
DRAM[1817] = 8'b1100101;
DRAM[1818] = 8'b1100101;
DRAM[1819] = 8'b1100110;
DRAM[1820] = 8'b1100110;
DRAM[1821] = 8'b1100111;
DRAM[1822] = 8'b1100111;
DRAM[1823] = 8'b1100111;
DRAM[1824] = 8'b1101000;
DRAM[1825] = 8'b1101000;
DRAM[1826] = 8'b1101001;
DRAM[1827] = 8'b1101010;
DRAM[1828] = 8'b1101100;
DRAM[1829] = 8'b1101101;
DRAM[1830] = 8'b1101110;
DRAM[1831] = 8'b1101111;
DRAM[1832] = 8'b1101101;
DRAM[1833] = 8'b1101101;
DRAM[1834] = 8'b1101110;
DRAM[1835] = 8'b1101111;
DRAM[1836] = 8'b1110000;
DRAM[1837] = 8'b1110000;
DRAM[1838] = 8'b1110001;
DRAM[1839] = 8'b1110010;
DRAM[1840] = 8'b1110000;
DRAM[1841] = 8'b1110000;
DRAM[1842] = 8'b1110000;
DRAM[1843] = 8'b1110000;
DRAM[1844] = 8'b1110000;
DRAM[1845] = 8'b1110000;
DRAM[1846] = 8'b1110000;
DRAM[1847] = 8'b1110000;
DRAM[1848] = 8'b1110001;
DRAM[1849] = 8'b1110001;
DRAM[1850] = 8'b1110001;
DRAM[1851] = 8'b1110001;
DRAM[1852] = 8'b1110001;
DRAM[1853] = 8'b1110001;
DRAM[1854] = 8'b1110001;
DRAM[1855] = 8'b1110001;
DRAM[1856] = 8'b1110000;
DRAM[1857] = 8'b1110000;
DRAM[1858] = 8'b1110000;
DRAM[1859] = 8'b1110001;
DRAM[1860] = 8'b1110001;
DRAM[1861] = 8'b1110010;
DRAM[1862] = 8'b1110010;
DRAM[1863] = 8'b1110011;
DRAM[1864] = 8'b1110000;
DRAM[1865] = 8'b1110001;
DRAM[1866] = 8'b1110001;
DRAM[1867] = 8'b1110001;
DRAM[1868] = 8'b1110001;
DRAM[1869] = 8'b1110000;
DRAM[1870] = 8'b1101111;
DRAM[1871] = 8'b1101110;
DRAM[1872] = 8'b1110000;
DRAM[1873] = 8'b1101111;
DRAM[1874] = 8'b1101110;
DRAM[1875] = 8'b1101101;
DRAM[1876] = 8'b1101101;
DRAM[1877] = 8'b1101101;
DRAM[1878] = 8'b1101110;
DRAM[1879] = 8'b1101110;
DRAM[1880] = 8'b1101110;
DRAM[1881] = 8'b1101110;
DRAM[1882] = 8'b1101110;
DRAM[1883] = 8'b1101110;
DRAM[1884] = 8'b1101110;
DRAM[1885] = 8'b1101110;
DRAM[1886] = 8'b1101110;
DRAM[1887] = 8'b1101110;
DRAM[1888] = 8'b1101111;
DRAM[1889] = 8'b1101111;
DRAM[1890] = 8'b1101110;
DRAM[1891] = 8'b1101110;
DRAM[1892] = 8'b1101111;
DRAM[1893] = 8'b1101111;
DRAM[1894] = 8'b1110000;
DRAM[1895] = 8'b1110001;
DRAM[1896] = 8'b1101111;
DRAM[1897] = 8'b1101111;
DRAM[1898] = 8'b1101111;
DRAM[1899] = 8'b1101110;
DRAM[1900] = 8'b1101110;
DRAM[1901] = 8'b1101110;
DRAM[1902] = 8'b1101101;
DRAM[1903] = 8'b1101101;
DRAM[1904] = 8'b1101101;
DRAM[1905] = 8'b1101101;
DRAM[1906] = 8'b1101101;
DRAM[1907] = 8'b1101101;
DRAM[1908] = 8'b1101101;
DRAM[1909] = 8'b1101101;
DRAM[1910] = 8'b1101101;
DRAM[1911] = 8'b1101101;
DRAM[1912] = 8'b1101100;
DRAM[1913] = 8'b1101100;
DRAM[1914] = 8'b1101100;
DRAM[1915] = 8'b1101100;
DRAM[1916] = 8'b1101100;
DRAM[1917] = 8'b1101100;
DRAM[1918] = 8'b1101100;
DRAM[1919] = 8'b1101100;
DRAM[1920] = 8'b1101111;
DRAM[1921] = 8'b1101110;
DRAM[1922] = 8'b1101110;
DRAM[1923] = 8'b1101101;
DRAM[1924] = 8'b1101101;
DRAM[1925] = 8'b1101100;
DRAM[1926] = 8'b1101100;
DRAM[1927] = 8'b1101100;
DRAM[1928] = 8'b1101011;
DRAM[1929] = 8'b1101100;
DRAM[1930] = 8'b1101101;
DRAM[1931] = 8'b1101110;
DRAM[1932] = 8'b1101110;
DRAM[1933] = 8'b1101110;
DRAM[1934] = 8'b1101110;
DRAM[1935] = 8'b1101101;
DRAM[1936] = 8'b1101101;
DRAM[1937] = 8'b1101110;
DRAM[1938] = 8'b1101111;
DRAM[1939] = 8'b1101111;
DRAM[1940] = 8'b1101111;
DRAM[1941] = 8'b1101111;
DRAM[1942] = 8'b1101110;
DRAM[1943] = 8'b1101101;
DRAM[1944] = 8'b1101100;
DRAM[1945] = 8'b1101100;
DRAM[1946] = 8'b1101100;
DRAM[1947] = 8'b1101100;
DRAM[1948] = 8'b1101100;
DRAM[1949] = 8'b1101100;
DRAM[1950] = 8'b1101100;
DRAM[1951] = 8'b1101100;
DRAM[1952] = 8'b1101010;
DRAM[1953] = 8'b1101011;
DRAM[1954] = 8'b1101011;
DRAM[1955] = 8'b1101010;
DRAM[1956] = 8'b1101001;
DRAM[1957] = 8'b1101000;
DRAM[1958] = 8'b1100111;
DRAM[1959] = 8'b1100110;
DRAM[1960] = 8'b1100101;
DRAM[1961] = 8'b1100101;
DRAM[1962] = 8'b1100110;
DRAM[1963] = 8'b1100111;
DRAM[1964] = 8'b1100110;
DRAM[1965] = 8'b1100101;
DRAM[1966] = 8'b1100100;
DRAM[1967] = 8'b1100010;
DRAM[1968] = 8'b1100011;
DRAM[1969] = 8'b1100011;
DRAM[1970] = 8'b1100011;
DRAM[1971] = 8'b1100010;
DRAM[1972] = 8'b1100010;
DRAM[1973] = 8'b1100010;
DRAM[1974] = 8'b1100001;
DRAM[1975] = 8'b1100001;
DRAM[1976] = 8'b1100001;
DRAM[1977] = 8'b1100001;
DRAM[1978] = 8'b1100000;
DRAM[1979] = 8'b1100000;
DRAM[1980] = 8'b1011111;
DRAM[1981] = 8'b1011110;
DRAM[1982] = 8'b1011101;
DRAM[1983] = 8'b1011101;
DRAM[1984] = 8'b1011100;
DRAM[1985] = 8'b1011011;
DRAM[1986] = 8'b1011010;
DRAM[1987] = 8'b1011010;
DRAM[1988] = 8'b1011001;
DRAM[1989] = 8'b1011000;
DRAM[1990] = 8'b1010111;
DRAM[1991] = 8'b1010111;
DRAM[1992] = 8'b1010111;
DRAM[1993] = 8'b1010111;
DRAM[1994] = 8'b1010111;
DRAM[1995] = 8'b1010110;
DRAM[1996] = 8'b1010110;
DRAM[1997] = 8'b1010110;
DRAM[1998] = 8'b1010101;
DRAM[1999] = 8'b1010101;
DRAM[2000] = 8'b1010010;
DRAM[2001] = 8'b1010010;
DRAM[2002] = 8'b1010010;
DRAM[2003] = 8'b1010001;
DRAM[2004] = 8'b1010001;
DRAM[2005] = 8'b1010000;
DRAM[2006] = 8'b1010000;
DRAM[2007] = 8'b1010000;
DRAM[2008] = 8'b1001110;
DRAM[2009] = 8'b1001110;
DRAM[2010] = 8'b1001111;
DRAM[2011] = 8'b1001111;
DRAM[2012] = 8'b1001111;
DRAM[2013] = 8'b1001110;
DRAM[2014] = 8'b1001101;
DRAM[2015] = 8'b1001101;
DRAM[2016] = 8'b1001011;
DRAM[2017] = 8'b1001011;
DRAM[2018] = 8'b1001011;
DRAM[2019] = 8'b1001010;
DRAM[2020] = 8'b1001010;
DRAM[2021] = 8'b1001010;
DRAM[2022] = 8'b1001001;
DRAM[2023] = 8'b1001001;
DRAM[2024] = 8'b1001000;
DRAM[2025] = 8'b1001000;
DRAM[2026] = 8'b1001000;
DRAM[2027] = 8'b1000111;
DRAM[2028] = 8'b1000111;
DRAM[2029] = 8'b1000110;
DRAM[2030] = 8'b1000110;
DRAM[2031] = 8'b1000110;
DRAM[2032] = 8'b1000100;
DRAM[2033] = 8'b1000100;
DRAM[2034] = 8'b1000100;
DRAM[2035] = 8'b1000011;
DRAM[2036] = 8'b1000011;
DRAM[2037] = 8'b1000010;
DRAM[2038] = 8'b1000010;
DRAM[2039] = 8'b1000010;
DRAM[2040] = 8'b1000010;
DRAM[2041] = 8'b1000010;
DRAM[2042] = 8'b1000010;
DRAM[2043] = 8'b1000001;
DRAM[2044] = 8'b1000001;
DRAM[2045] = 8'b1000001;
DRAM[2046] = 8'b1000000;
DRAM[2047] = 8'b1000000;
DRAM[2048] = 8'b1011010;
DRAM[2049] = 8'b1011011;
DRAM[2050] = 8'b1011100;
DRAM[2051] = 8'b1011101;
DRAM[2052] = 8'b1011111;
DRAM[2053] = 8'b1100000;
DRAM[2054] = 8'b1100001;
DRAM[2055] = 8'b1100001;
DRAM[2056] = 8'b1100000;
DRAM[2057] = 8'b1100001;
DRAM[2058] = 8'b1100010;
DRAM[2059] = 8'b1100010;
DRAM[2060] = 8'b1100011;
DRAM[2061] = 8'b1100100;
DRAM[2062] = 8'b1100101;
DRAM[2063] = 8'b1100101;
DRAM[2064] = 8'b1100100;
DRAM[2065] = 8'b1100100;
DRAM[2066] = 8'b1100101;
DRAM[2067] = 8'b1100110;
DRAM[2068] = 8'b1100110;
DRAM[2069] = 8'b1100111;
DRAM[2070] = 8'b1101000;
DRAM[2071] = 8'b1101000;
DRAM[2072] = 8'b1100110;
DRAM[2073] = 8'b1100111;
DRAM[2074] = 8'b1101000;
DRAM[2075] = 8'b1101001;
DRAM[2076] = 8'b1101001;
DRAM[2077] = 8'b1101001;
DRAM[2078] = 8'b1101001;
DRAM[2079] = 8'b1101000;
DRAM[2080] = 8'b1101010;
DRAM[2081] = 8'b1101010;
DRAM[2082] = 8'b1101010;
DRAM[2083] = 8'b1101011;
DRAM[2084] = 8'b1101011;
DRAM[2085] = 8'b1101100;
DRAM[2086] = 8'b1101100;
DRAM[2087] = 8'b1101100;
DRAM[2088] = 8'b1101100;
DRAM[2089] = 8'b1101100;
DRAM[2090] = 8'b1101100;
DRAM[2091] = 8'b1101101;
DRAM[2092] = 8'b1101101;
DRAM[2093] = 8'b1101110;
DRAM[2094] = 8'b1101110;
DRAM[2095] = 8'b1101110;
DRAM[2096] = 8'b1110010;
DRAM[2097] = 8'b1110001;
DRAM[2098] = 8'b1110000;
DRAM[2099] = 8'b1101111;
DRAM[2100] = 8'b1110000;
DRAM[2101] = 8'b1110001;
DRAM[2102] = 8'b1110011;
DRAM[2103] = 8'b1110100;
DRAM[2104] = 8'b1110001;
DRAM[2105] = 8'b1110001;
DRAM[2106] = 8'b1110001;
DRAM[2107] = 8'b1110001;
DRAM[2108] = 8'b1110001;
DRAM[2109] = 8'b1110001;
DRAM[2110] = 8'b1110001;
DRAM[2111] = 8'b1110001;
DRAM[2112] = 8'b1110010;
DRAM[2113] = 8'b1110010;
DRAM[2114] = 8'b1110010;
DRAM[2115] = 8'b1110010;
DRAM[2116] = 8'b1110010;
DRAM[2117] = 8'b1110010;
DRAM[2118] = 8'b1110010;
DRAM[2119] = 8'b1110010;
DRAM[2120] = 8'b1110001;
DRAM[2121] = 8'b1110001;
DRAM[2122] = 8'b1110001;
DRAM[2123] = 8'b1110001;
DRAM[2124] = 8'b1110001;
DRAM[2125] = 8'b1110001;
DRAM[2126] = 8'b1110001;
DRAM[2127] = 8'b1110001;
DRAM[2128] = 8'b1110011;
DRAM[2129] = 8'b1110010;
DRAM[2130] = 8'b1110001;
DRAM[2131] = 8'b1110000;
DRAM[2132] = 8'b1101111;
DRAM[2133] = 8'b1101110;
DRAM[2134] = 8'b1101110;
DRAM[2135] = 8'b1101101;
DRAM[2136] = 8'b1101111;
DRAM[2137] = 8'b1101111;
DRAM[2138] = 8'b1101111;
DRAM[2139] = 8'b1101111;
DRAM[2140] = 8'b1101111;
DRAM[2141] = 8'b1101111;
DRAM[2142] = 8'b1101111;
DRAM[2143] = 8'b1101111;
DRAM[2144] = 8'b1110001;
DRAM[2145] = 8'b1110000;
DRAM[2146] = 8'b1101111;
DRAM[2147] = 8'b1101111;
DRAM[2148] = 8'b1110001;
DRAM[2149] = 8'b1110001;
DRAM[2150] = 8'b1110000;
DRAM[2151] = 8'b1101111;
DRAM[2152] = 8'b1110000;
DRAM[2153] = 8'b1110001;
DRAM[2154] = 8'b1110001;
DRAM[2155] = 8'b1110010;
DRAM[2156] = 8'b1110010;
DRAM[2157] = 8'b1110001;
DRAM[2158] = 8'b1110001;
DRAM[2159] = 8'b1110000;
DRAM[2160] = 8'b1101101;
DRAM[2161] = 8'b1101101;
DRAM[2162] = 8'b1101101;
DRAM[2163] = 8'b1101101;
DRAM[2164] = 8'b1101101;
DRAM[2165] = 8'b1101101;
DRAM[2166] = 8'b1101101;
DRAM[2167] = 8'b1101101;
DRAM[2168] = 8'b1101101;
DRAM[2169] = 8'b1101101;
DRAM[2170] = 8'b1101101;
DRAM[2171] = 8'b1101101;
DRAM[2172] = 8'b1101101;
DRAM[2173] = 8'b1101101;
DRAM[2174] = 8'b1101101;
DRAM[2175] = 8'b1101101;
DRAM[2176] = 8'b1101101;
DRAM[2177] = 8'b1101101;
DRAM[2178] = 8'b1101101;
DRAM[2179] = 8'b1101101;
DRAM[2180] = 8'b1101101;
DRAM[2181] = 8'b1101101;
DRAM[2182] = 8'b1101101;
DRAM[2183] = 8'b1101101;
DRAM[2184] = 8'b1101100;
DRAM[2185] = 8'b1101101;
DRAM[2186] = 8'b1101101;
DRAM[2187] = 8'b1101110;
DRAM[2188] = 8'b1101110;
DRAM[2189] = 8'b1101101;
DRAM[2190] = 8'b1101101;
DRAM[2191] = 8'b1101100;
DRAM[2192] = 8'b1101110;
DRAM[2193] = 8'b1101111;
DRAM[2194] = 8'b1101111;
DRAM[2195] = 8'b1110000;
DRAM[2196] = 8'b1110000;
DRAM[2197] = 8'b1101111;
DRAM[2198] = 8'b1101111;
DRAM[2199] = 8'b1101110;
DRAM[2200] = 8'b1101100;
DRAM[2201] = 8'b1101100;
DRAM[2202] = 8'b1101100;
DRAM[2203] = 8'b1101100;
DRAM[2204] = 8'b1101100;
DRAM[2205] = 8'b1101100;
DRAM[2206] = 8'b1101100;
DRAM[2207] = 8'b1101100;
DRAM[2208] = 8'b1101010;
DRAM[2209] = 8'b1101010;
DRAM[2210] = 8'b1101010;
DRAM[2211] = 8'b1101010;
DRAM[2212] = 8'b1101010;
DRAM[2213] = 8'b1101010;
DRAM[2214] = 8'b1101010;
DRAM[2215] = 8'b1101010;
DRAM[2216] = 8'b1100111;
DRAM[2217] = 8'b1100111;
DRAM[2218] = 8'b1100110;
DRAM[2219] = 8'b1100110;
DRAM[2220] = 8'b1100110;
DRAM[2221] = 8'b1100101;
DRAM[2222] = 8'b1100101;
DRAM[2223] = 8'b1100101;
DRAM[2224] = 8'b1100110;
DRAM[2225] = 8'b1100110;
DRAM[2226] = 8'b1100101;
DRAM[2227] = 8'b1100100;
DRAM[2228] = 8'b1100011;
DRAM[2229] = 8'b1100011;
DRAM[2230] = 8'b1100010;
DRAM[2231] = 8'b1100010;
DRAM[2232] = 8'b1100001;
DRAM[2233] = 8'b1100001;
DRAM[2234] = 8'b1100000;
DRAM[2235] = 8'b1011111;
DRAM[2236] = 8'b1011110;
DRAM[2237] = 8'b1011110;
DRAM[2238] = 8'b1011101;
DRAM[2239] = 8'b1011101;
DRAM[2240] = 8'b1011100;
DRAM[2241] = 8'b1011100;
DRAM[2242] = 8'b1011011;
DRAM[2243] = 8'b1011010;
DRAM[2244] = 8'b1011001;
DRAM[2245] = 8'b1011001;
DRAM[2246] = 8'b1011000;
DRAM[2247] = 8'b1011000;
DRAM[2248] = 8'b1011011;
DRAM[2249] = 8'b1011010;
DRAM[2250] = 8'b1011001;
DRAM[2251] = 8'b1011000;
DRAM[2252] = 8'b1010110;
DRAM[2253] = 8'b1010101;
DRAM[2254] = 8'b1010100;
DRAM[2255] = 8'b1010011;
DRAM[2256] = 8'b1010101;
DRAM[2257] = 8'b1010100;
DRAM[2258] = 8'b1010011;
DRAM[2259] = 8'b1010010;
DRAM[2260] = 8'b1010001;
DRAM[2261] = 8'b1010000;
DRAM[2262] = 8'b1010001;
DRAM[2263] = 8'b1010001;
DRAM[2264] = 8'b1001111;
DRAM[2265] = 8'b1001111;
DRAM[2266] = 8'b1001111;
DRAM[2267] = 8'b1001111;
DRAM[2268] = 8'b1001111;
DRAM[2269] = 8'b1001111;
DRAM[2270] = 8'b1001111;
DRAM[2271] = 8'b1001111;
DRAM[2272] = 8'b1001101;
DRAM[2273] = 8'b1001100;
DRAM[2274] = 8'b1001011;
DRAM[2275] = 8'b1001010;
DRAM[2276] = 8'b1001010;
DRAM[2277] = 8'b1001010;
DRAM[2278] = 8'b1001010;
DRAM[2279] = 8'b1001011;
DRAM[2280] = 8'b1001001;
DRAM[2281] = 8'b1001001;
DRAM[2282] = 8'b1001000;
DRAM[2283] = 8'b1000111;
DRAM[2284] = 8'b1000110;
DRAM[2285] = 8'b1000110;
DRAM[2286] = 8'b1000101;
DRAM[2287] = 8'b1000100;
DRAM[2288] = 8'b1000101;
DRAM[2289] = 8'b1000101;
DRAM[2290] = 8'b1000100;
DRAM[2291] = 8'b1000100;
DRAM[2292] = 8'b1000100;
DRAM[2293] = 8'b1000011;
DRAM[2294] = 8'b1000011;
DRAM[2295] = 8'b1000011;
DRAM[2296] = 8'b1000010;
DRAM[2297] = 8'b1000010;
DRAM[2298] = 8'b1000010;
DRAM[2299] = 8'b1000001;
DRAM[2300] = 8'b1000001;
DRAM[2301] = 8'b1000000;
DRAM[2302] = 8'b1000000;
DRAM[2303] = 8'b1000000;
DRAM[2304] = 8'b1011011;
DRAM[2305] = 8'b1011011;
DRAM[2306] = 8'b1011100;
DRAM[2307] = 8'b1011110;
DRAM[2308] = 8'b1011111;
DRAM[2309] = 8'b1100000;
DRAM[2310] = 8'b1100001;
DRAM[2311] = 8'b1100010;
DRAM[2312] = 8'b1100010;
DRAM[2313] = 8'b1100010;
DRAM[2314] = 8'b1100011;
DRAM[2315] = 8'b1100100;
DRAM[2316] = 8'b1100101;
DRAM[2317] = 8'b1100110;
DRAM[2318] = 8'b1100110;
DRAM[2319] = 8'b1100111;
DRAM[2320] = 8'b1100011;
DRAM[2321] = 8'b1100011;
DRAM[2322] = 8'b1100100;
DRAM[2323] = 8'b1100100;
DRAM[2324] = 8'b1100101;
DRAM[2325] = 8'b1100110;
DRAM[2326] = 8'b1100111;
DRAM[2327] = 8'b1100111;
DRAM[2328] = 8'b1100110;
DRAM[2329] = 8'b1100110;
DRAM[2330] = 8'b1100111;
DRAM[2331] = 8'b1101000;
DRAM[2332] = 8'b1101001;
DRAM[2333] = 8'b1101001;
DRAM[2334] = 8'b1101000;
DRAM[2335] = 8'b1101000;
DRAM[2336] = 8'b1101011;
DRAM[2337] = 8'b1101011;
DRAM[2338] = 8'b1101100;
DRAM[2339] = 8'b1101100;
DRAM[2340] = 8'b1101101;
DRAM[2341] = 8'b1101101;
DRAM[2342] = 8'b1101101;
DRAM[2343] = 8'b1101101;
DRAM[2344] = 8'b1101100;
DRAM[2345] = 8'b1101100;
DRAM[2346] = 8'b1101101;
DRAM[2347] = 8'b1101101;
DRAM[2348] = 8'b1101101;
DRAM[2349] = 8'b1101110;
DRAM[2350] = 8'b1101110;
DRAM[2351] = 8'b1101110;
DRAM[2352] = 8'b1110001;
DRAM[2353] = 8'b1110001;
DRAM[2354] = 8'b1110000;
DRAM[2355] = 8'b1110000;
DRAM[2356] = 8'b1110000;
DRAM[2357] = 8'b1110001;
DRAM[2358] = 8'b1110011;
DRAM[2359] = 8'b1110100;
DRAM[2360] = 8'b1110010;
DRAM[2361] = 8'b1110010;
DRAM[2362] = 8'b1110010;
DRAM[2363] = 8'b1110010;
DRAM[2364] = 8'b1110010;
DRAM[2365] = 8'b1110010;
DRAM[2366] = 8'b1110010;
DRAM[2367] = 8'b1110010;
DRAM[2368] = 8'b1110010;
DRAM[2369] = 8'b1110010;
DRAM[2370] = 8'b1110010;
DRAM[2371] = 8'b1110010;
DRAM[2372] = 8'b1110010;
DRAM[2373] = 8'b1110010;
DRAM[2374] = 8'b1110010;
DRAM[2375] = 8'b1110010;
DRAM[2376] = 8'b1110001;
DRAM[2377] = 8'b1110001;
DRAM[2378] = 8'b1110001;
DRAM[2379] = 8'b1110001;
DRAM[2380] = 8'b1110001;
DRAM[2381] = 8'b1110001;
DRAM[2382] = 8'b1110001;
DRAM[2383] = 8'b1110001;
DRAM[2384] = 8'b1110010;
DRAM[2385] = 8'b1110010;
DRAM[2386] = 8'b1110001;
DRAM[2387] = 8'b1110001;
DRAM[2388] = 8'b1110000;
DRAM[2389] = 8'b1101111;
DRAM[2390] = 8'b1101111;
DRAM[2391] = 8'b1101111;
DRAM[2392] = 8'b1101111;
DRAM[2393] = 8'b1101111;
DRAM[2394] = 8'b1101111;
DRAM[2395] = 8'b1101111;
DRAM[2396] = 8'b1101111;
DRAM[2397] = 8'b1101111;
DRAM[2398] = 8'b1101111;
DRAM[2399] = 8'b1101111;
DRAM[2400] = 8'b1110001;
DRAM[2401] = 8'b1110000;
DRAM[2402] = 8'b1101111;
DRAM[2403] = 8'b1101111;
DRAM[2404] = 8'b1110001;
DRAM[2405] = 8'b1110010;
DRAM[2406] = 8'b1110000;
DRAM[2407] = 8'b1101111;
DRAM[2408] = 8'b1110000;
DRAM[2409] = 8'b1110000;
DRAM[2410] = 8'b1110001;
DRAM[2411] = 8'b1110001;
DRAM[2412] = 8'b1110001;
DRAM[2413] = 8'b1110001;
DRAM[2414] = 8'b1110000;
DRAM[2415] = 8'b1110000;
DRAM[2416] = 8'b1101101;
DRAM[2417] = 8'b1101101;
DRAM[2418] = 8'b1101101;
DRAM[2419] = 8'b1101101;
DRAM[2420] = 8'b1101101;
DRAM[2421] = 8'b1101101;
DRAM[2422] = 8'b1101101;
DRAM[2423] = 8'b1101101;
DRAM[2424] = 8'b1101101;
DRAM[2425] = 8'b1101101;
DRAM[2426] = 8'b1101101;
DRAM[2427] = 8'b1101101;
DRAM[2428] = 8'b1101101;
DRAM[2429] = 8'b1101101;
DRAM[2430] = 8'b1101101;
DRAM[2431] = 8'b1101101;
DRAM[2432] = 8'b1101101;
DRAM[2433] = 8'b1101101;
DRAM[2434] = 8'b1101101;
DRAM[2435] = 8'b1101101;
DRAM[2436] = 8'b1101101;
DRAM[2437] = 8'b1101101;
DRAM[2438] = 8'b1101101;
DRAM[2439] = 8'b1101101;
DRAM[2440] = 8'b1101110;
DRAM[2441] = 8'b1101110;
DRAM[2442] = 8'b1101111;
DRAM[2443] = 8'b1101111;
DRAM[2444] = 8'b1101111;
DRAM[2445] = 8'b1101111;
DRAM[2446] = 8'b1101110;
DRAM[2447] = 8'b1101110;
DRAM[2448] = 8'b1101110;
DRAM[2449] = 8'b1101110;
DRAM[2450] = 8'b1101111;
DRAM[2451] = 8'b1110000;
DRAM[2452] = 8'b1110000;
DRAM[2453] = 8'b1101111;
DRAM[2454] = 8'b1101110;
DRAM[2455] = 8'b1101110;
DRAM[2456] = 8'b1101100;
DRAM[2457] = 8'b1101100;
DRAM[2458] = 8'b1101100;
DRAM[2459] = 8'b1101100;
DRAM[2460] = 8'b1101100;
DRAM[2461] = 8'b1101100;
DRAM[2462] = 8'b1101100;
DRAM[2463] = 8'b1101100;
DRAM[2464] = 8'b1101010;
DRAM[2465] = 8'b1101010;
DRAM[2466] = 8'b1101010;
DRAM[2467] = 8'b1101010;
DRAM[2468] = 8'b1101010;
DRAM[2469] = 8'b1101010;
DRAM[2470] = 8'b1101010;
DRAM[2471] = 8'b1101010;
DRAM[2472] = 8'b1101000;
DRAM[2473] = 8'b1101000;
DRAM[2474] = 8'b1100111;
DRAM[2475] = 8'b1100111;
DRAM[2476] = 8'b1100111;
DRAM[2477] = 8'b1100110;
DRAM[2478] = 8'b1100110;
DRAM[2479] = 8'b1100110;
DRAM[2480] = 8'b1100110;
DRAM[2481] = 8'b1100110;
DRAM[2482] = 8'b1100101;
DRAM[2483] = 8'b1100101;
DRAM[2484] = 8'b1100100;
DRAM[2485] = 8'b1100011;
DRAM[2486] = 8'b1100010;
DRAM[2487] = 8'b1100010;
DRAM[2488] = 8'b1100001;
DRAM[2489] = 8'b1100001;
DRAM[2490] = 8'b1100000;
DRAM[2491] = 8'b1100000;
DRAM[2492] = 8'b1011111;
DRAM[2493] = 8'b1011110;
DRAM[2494] = 8'b1011101;
DRAM[2495] = 8'b1011101;
DRAM[2496] = 8'b1011100;
DRAM[2497] = 8'b1011100;
DRAM[2498] = 8'b1011011;
DRAM[2499] = 8'b1011011;
DRAM[2500] = 8'b1011010;
DRAM[2501] = 8'b1011001;
DRAM[2502] = 8'b1011000;
DRAM[2503] = 8'b1011000;
DRAM[2504] = 8'b1011010;
DRAM[2505] = 8'b1011001;
DRAM[2506] = 8'b1011001;
DRAM[2507] = 8'b1011000;
DRAM[2508] = 8'b1010111;
DRAM[2509] = 8'b1010110;
DRAM[2510] = 8'b1010101;
DRAM[2511] = 8'b1010100;
DRAM[2512] = 8'b1010101;
DRAM[2513] = 8'b1010100;
DRAM[2514] = 8'b1010011;
DRAM[2515] = 8'b1010010;
DRAM[2516] = 8'b1010001;
DRAM[2517] = 8'b1010001;
DRAM[2518] = 8'b1010001;
DRAM[2519] = 8'b1010001;
DRAM[2520] = 8'b1001111;
DRAM[2521] = 8'b1001111;
DRAM[2522] = 8'b1001111;
DRAM[2523] = 8'b1001111;
DRAM[2524] = 8'b1001111;
DRAM[2525] = 8'b1001111;
DRAM[2526] = 8'b1001111;
DRAM[2527] = 8'b1001111;
DRAM[2528] = 8'b1001101;
DRAM[2529] = 8'b1001100;
DRAM[2530] = 8'b1001011;
DRAM[2531] = 8'b1001011;
DRAM[2532] = 8'b1001010;
DRAM[2533] = 8'b1001010;
DRAM[2534] = 8'b1001011;
DRAM[2535] = 8'b1001011;
DRAM[2536] = 8'b1001010;
DRAM[2537] = 8'b1001001;
DRAM[2538] = 8'b1001001;
DRAM[2539] = 8'b1001000;
DRAM[2540] = 8'b1000111;
DRAM[2541] = 8'b1000110;
DRAM[2542] = 8'b1000101;
DRAM[2543] = 8'b1000101;
DRAM[2544] = 8'b1000101;
DRAM[2545] = 8'b1000101;
DRAM[2546] = 8'b1000101;
DRAM[2547] = 8'b1000100;
DRAM[2548] = 8'b1000100;
DRAM[2549] = 8'b1000100;
DRAM[2550] = 8'b1000011;
DRAM[2551] = 8'b1000011;
DRAM[2552] = 8'b1000010;
DRAM[2553] = 8'b1000010;
DRAM[2554] = 8'b1000010;
DRAM[2555] = 8'b1000001;
DRAM[2556] = 8'b1000001;
DRAM[2557] = 8'b1000001;
DRAM[2558] = 8'b1000000;
DRAM[2559] = 8'b1000000;
DRAM[2560] = 8'b1011100;
DRAM[2561] = 8'b1011100;
DRAM[2562] = 8'b1011101;
DRAM[2563] = 8'b1011110;
DRAM[2564] = 8'b1011111;
DRAM[2565] = 8'b1100000;
DRAM[2566] = 8'b1100001;
DRAM[2567] = 8'b1100010;
DRAM[2568] = 8'b1100011;
DRAM[2569] = 8'b1100100;
DRAM[2570] = 8'b1100100;
DRAM[2571] = 8'b1100101;
DRAM[2572] = 8'b1100110;
DRAM[2573] = 8'b1100110;
DRAM[2574] = 8'b1100111;
DRAM[2575] = 8'b1100111;
DRAM[2576] = 8'b1100010;
DRAM[2577] = 8'b1100010;
DRAM[2578] = 8'b1100011;
DRAM[2579] = 8'b1100100;
DRAM[2580] = 8'b1100101;
DRAM[2581] = 8'b1100101;
DRAM[2582] = 8'b1100110;
DRAM[2583] = 8'b1100110;
DRAM[2584] = 8'b1100101;
DRAM[2585] = 8'b1100110;
DRAM[2586] = 8'b1100111;
DRAM[2587] = 8'b1101000;
DRAM[2588] = 8'b1101000;
DRAM[2589] = 8'b1101000;
DRAM[2590] = 8'b1101000;
DRAM[2591] = 8'b1101000;
DRAM[2592] = 8'b1101101;
DRAM[2593] = 8'b1101101;
DRAM[2594] = 8'b1101101;
DRAM[2595] = 8'b1101101;
DRAM[2596] = 8'b1101110;
DRAM[2597] = 8'b1101110;
DRAM[2598] = 8'b1101111;
DRAM[2599] = 8'b1101111;
DRAM[2600] = 8'b1101100;
DRAM[2601] = 8'b1101101;
DRAM[2602] = 8'b1101101;
DRAM[2603] = 8'b1101101;
DRAM[2604] = 8'b1101110;
DRAM[2605] = 8'b1101110;
DRAM[2606] = 8'b1101110;
DRAM[2607] = 8'b1101110;
DRAM[2608] = 8'b1110001;
DRAM[2609] = 8'b1110001;
DRAM[2610] = 8'b1110000;
DRAM[2611] = 8'b1110000;
DRAM[2612] = 8'b1110001;
DRAM[2613] = 8'b1110010;
DRAM[2614] = 8'b1110011;
DRAM[2615] = 8'b1110011;
DRAM[2616] = 8'b1110011;
DRAM[2617] = 8'b1110011;
DRAM[2618] = 8'b1110011;
DRAM[2619] = 8'b1110011;
DRAM[2620] = 8'b1110011;
DRAM[2621] = 8'b1110011;
DRAM[2622] = 8'b1110011;
DRAM[2623] = 8'b1110011;
DRAM[2624] = 8'b1110010;
DRAM[2625] = 8'b1110010;
DRAM[2626] = 8'b1110010;
DRAM[2627] = 8'b1110010;
DRAM[2628] = 8'b1110010;
DRAM[2629] = 8'b1110010;
DRAM[2630] = 8'b1110010;
DRAM[2631] = 8'b1110010;
DRAM[2632] = 8'b1110001;
DRAM[2633] = 8'b1110001;
DRAM[2634] = 8'b1110001;
DRAM[2635] = 8'b1110001;
DRAM[2636] = 8'b1110001;
DRAM[2637] = 8'b1110001;
DRAM[2638] = 8'b1110001;
DRAM[2639] = 8'b1110001;
DRAM[2640] = 8'b1110001;
DRAM[2641] = 8'b1110001;
DRAM[2642] = 8'b1110001;
DRAM[2643] = 8'b1110001;
DRAM[2644] = 8'b1110001;
DRAM[2645] = 8'b1110001;
DRAM[2646] = 8'b1110000;
DRAM[2647] = 8'b1110000;
DRAM[2648] = 8'b1101111;
DRAM[2649] = 8'b1101111;
DRAM[2650] = 8'b1101111;
DRAM[2651] = 8'b1101111;
DRAM[2652] = 8'b1101111;
DRAM[2653] = 8'b1101111;
DRAM[2654] = 8'b1101111;
DRAM[2655] = 8'b1101111;
DRAM[2656] = 8'b1110010;
DRAM[2657] = 8'b1110000;
DRAM[2658] = 8'b1101111;
DRAM[2659] = 8'b1110000;
DRAM[2660] = 8'b1110001;
DRAM[2661] = 8'b1110010;
DRAM[2662] = 8'b1110001;
DRAM[2663] = 8'b1101111;
DRAM[2664] = 8'b1101111;
DRAM[2665] = 8'b1110000;
DRAM[2666] = 8'b1110000;
DRAM[2667] = 8'b1110001;
DRAM[2668] = 8'b1110001;
DRAM[2669] = 8'b1110000;
DRAM[2670] = 8'b1110000;
DRAM[2671] = 8'b1101111;
DRAM[2672] = 8'b1101110;
DRAM[2673] = 8'b1101110;
DRAM[2674] = 8'b1101110;
DRAM[2675] = 8'b1101110;
DRAM[2676] = 8'b1101110;
DRAM[2677] = 8'b1101110;
DRAM[2678] = 8'b1101110;
DRAM[2679] = 8'b1101110;
DRAM[2680] = 8'b1101110;
DRAM[2681] = 8'b1101110;
DRAM[2682] = 8'b1101110;
DRAM[2683] = 8'b1101110;
DRAM[2684] = 8'b1101110;
DRAM[2685] = 8'b1101110;
DRAM[2686] = 8'b1101110;
DRAM[2687] = 8'b1101110;
DRAM[2688] = 8'b1101110;
DRAM[2689] = 8'b1101110;
DRAM[2690] = 8'b1101110;
DRAM[2691] = 8'b1101110;
DRAM[2692] = 8'b1101110;
DRAM[2693] = 8'b1101110;
DRAM[2694] = 8'b1101110;
DRAM[2695] = 8'b1101110;
DRAM[2696] = 8'b1101111;
DRAM[2697] = 8'b1110000;
DRAM[2698] = 8'b1110000;
DRAM[2699] = 8'b1110001;
DRAM[2700] = 8'b1110001;
DRAM[2701] = 8'b1110000;
DRAM[2702] = 8'b1110000;
DRAM[2703] = 8'b1101111;
DRAM[2704] = 8'b1101110;
DRAM[2705] = 8'b1101110;
DRAM[2706] = 8'b1101111;
DRAM[2707] = 8'b1101111;
DRAM[2708] = 8'b1101111;
DRAM[2709] = 8'b1101111;
DRAM[2710] = 8'b1101110;
DRAM[2711] = 8'b1101110;
DRAM[2712] = 8'b1101101;
DRAM[2713] = 8'b1101101;
DRAM[2714] = 8'b1101101;
DRAM[2715] = 8'b1101101;
DRAM[2716] = 8'b1101101;
DRAM[2717] = 8'b1101101;
DRAM[2718] = 8'b1101101;
DRAM[2719] = 8'b1101101;
DRAM[2720] = 8'b1101011;
DRAM[2721] = 8'b1101011;
DRAM[2722] = 8'b1101011;
DRAM[2723] = 8'b1101011;
DRAM[2724] = 8'b1101011;
DRAM[2725] = 8'b1101011;
DRAM[2726] = 8'b1101011;
DRAM[2727] = 8'b1101011;
DRAM[2728] = 8'b1101001;
DRAM[2729] = 8'b1101001;
DRAM[2730] = 8'b1101001;
DRAM[2731] = 8'b1101000;
DRAM[2732] = 8'b1101000;
DRAM[2733] = 8'b1101000;
DRAM[2734] = 8'b1100111;
DRAM[2735] = 8'b1100111;
DRAM[2736] = 8'b1100111;
DRAM[2737] = 8'b1100111;
DRAM[2738] = 8'b1100110;
DRAM[2739] = 8'b1100101;
DRAM[2740] = 8'b1100100;
DRAM[2741] = 8'b1100100;
DRAM[2742] = 8'b1100011;
DRAM[2743] = 8'b1100011;
DRAM[2744] = 8'b1100010;
DRAM[2745] = 8'b1100010;
DRAM[2746] = 8'b1100001;
DRAM[2747] = 8'b1100000;
DRAM[2748] = 8'b1011111;
DRAM[2749] = 8'b1011111;
DRAM[2750] = 8'b1011110;
DRAM[2751] = 8'b1011110;
DRAM[2752] = 8'b1011101;
DRAM[2753] = 8'b1011101;
DRAM[2754] = 8'b1011100;
DRAM[2755] = 8'b1011011;
DRAM[2756] = 8'b1011010;
DRAM[2757] = 8'b1011010;
DRAM[2758] = 8'b1011001;
DRAM[2759] = 8'b1011001;
DRAM[2760] = 8'b1011001;
DRAM[2761] = 8'b1011001;
DRAM[2762] = 8'b1011000;
DRAM[2763] = 8'b1011000;
DRAM[2764] = 8'b1010111;
DRAM[2765] = 8'b1010111;
DRAM[2766] = 8'b1010110;
DRAM[2767] = 8'b1010110;
DRAM[2768] = 8'b1010101;
DRAM[2769] = 8'b1010101;
DRAM[2770] = 8'b1010011;
DRAM[2771] = 8'b1010010;
DRAM[2772] = 8'b1010001;
DRAM[2773] = 8'b1010001;
DRAM[2774] = 8'b1010001;
DRAM[2775] = 8'b1010001;
DRAM[2776] = 8'b1001111;
DRAM[2777] = 8'b1001111;
DRAM[2778] = 8'b1001111;
DRAM[2779] = 8'b1001111;
DRAM[2780] = 8'b1001111;
DRAM[2781] = 8'b1001111;
DRAM[2782] = 8'b1001111;
DRAM[2783] = 8'b1001111;
DRAM[2784] = 8'b1001101;
DRAM[2785] = 8'b1001101;
DRAM[2786] = 8'b1001100;
DRAM[2787] = 8'b1001011;
DRAM[2788] = 8'b1001010;
DRAM[2789] = 8'b1001010;
DRAM[2790] = 8'b1001011;
DRAM[2791] = 8'b1001011;
DRAM[2792] = 8'b1001010;
DRAM[2793] = 8'b1001001;
DRAM[2794] = 8'b1001001;
DRAM[2795] = 8'b1001000;
DRAM[2796] = 8'b1000111;
DRAM[2797] = 8'b1000111;
DRAM[2798] = 8'b1000110;
DRAM[2799] = 8'b1000110;
DRAM[2800] = 8'b1000110;
DRAM[2801] = 8'b1000110;
DRAM[2802] = 8'b1000101;
DRAM[2803] = 8'b1000101;
DRAM[2804] = 8'b1000101;
DRAM[2805] = 8'b1000100;
DRAM[2806] = 8'b1000100;
DRAM[2807] = 8'b1000100;
DRAM[2808] = 8'b1000010;
DRAM[2809] = 8'b1000010;
DRAM[2810] = 8'b1000010;
DRAM[2811] = 8'b1000010;
DRAM[2812] = 8'b1000001;
DRAM[2813] = 8'b1000001;
DRAM[2814] = 8'b1000001;
DRAM[2815] = 8'b1000000;
DRAM[2816] = 8'b1011101;
DRAM[2817] = 8'b1011110;
DRAM[2818] = 8'b1011110;
DRAM[2819] = 8'b1011111;
DRAM[2820] = 8'b1100000;
DRAM[2821] = 8'b1100001;
DRAM[2822] = 8'b1100010;
DRAM[2823] = 8'b1100010;
DRAM[2824] = 8'b1100011;
DRAM[2825] = 8'b1100100;
DRAM[2826] = 8'b1100100;
DRAM[2827] = 8'b1100100;
DRAM[2828] = 8'b1100101;
DRAM[2829] = 8'b1100101;
DRAM[2830] = 8'b1100110;
DRAM[2831] = 8'b1100110;
DRAM[2832] = 8'b1100011;
DRAM[2833] = 8'b1100011;
DRAM[2834] = 8'b1100100;
DRAM[2835] = 8'b1100101;
DRAM[2836] = 8'b1100110;
DRAM[2837] = 8'b1100110;
DRAM[2838] = 8'b1100111;
DRAM[2839] = 8'b1100111;
DRAM[2840] = 8'b1100110;
DRAM[2841] = 8'b1100110;
DRAM[2842] = 8'b1100111;
DRAM[2843] = 8'b1101000;
DRAM[2844] = 8'b1101000;
DRAM[2845] = 8'b1101000;
DRAM[2846] = 8'b1101000;
DRAM[2847] = 8'b1101000;
DRAM[2848] = 8'b1101100;
DRAM[2849] = 8'b1101101;
DRAM[2850] = 8'b1101101;
DRAM[2851] = 8'b1101101;
DRAM[2852] = 8'b1101110;
DRAM[2853] = 8'b1101110;
DRAM[2854] = 8'b1101110;
DRAM[2855] = 8'b1101111;
DRAM[2856] = 8'b1101101;
DRAM[2857] = 8'b1101101;
DRAM[2858] = 8'b1101101;
DRAM[2859] = 8'b1101110;
DRAM[2860] = 8'b1101110;
DRAM[2861] = 8'b1101110;
DRAM[2862] = 8'b1101111;
DRAM[2863] = 8'b1101111;
DRAM[2864] = 8'b1110001;
DRAM[2865] = 8'b1110001;
DRAM[2866] = 8'b1110001;
DRAM[2867] = 8'b1110001;
DRAM[2868] = 8'b1110010;
DRAM[2869] = 8'b1110010;
DRAM[2870] = 8'b1110011;
DRAM[2871] = 8'b1110011;
DRAM[2872] = 8'b1110100;
DRAM[2873] = 8'b1110100;
DRAM[2874] = 8'b1110100;
DRAM[2875] = 8'b1110100;
DRAM[2876] = 8'b1110100;
DRAM[2877] = 8'b1110100;
DRAM[2878] = 8'b1110100;
DRAM[2879] = 8'b1110100;
DRAM[2880] = 8'b1110011;
DRAM[2881] = 8'b1110011;
DRAM[2882] = 8'b1110011;
DRAM[2883] = 8'b1110011;
DRAM[2884] = 8'b1110011;
DRAM[2885] = 8'b1110011;
DRAM[2886] = 8'b1110011;
DRAM[2887] = 8'b1110011;
DRAM[2888] = 8'b1110010;
DRAM[2889] = 8'b1110010;
DRAM[2890] = 8'b1110010;
DRAM[2891] = 8'b1110010;
DRAM[2892] = 8'b1110010;
DRAM[2893] = 8'b1110010;
DRAM[2894] = 8'b1110010;
DRAM[2895] = 8'b1110010;
DRAM[2896] = 8'b1110001;
DRAM[2897] = 8'b1110001;
DRAM[2898] = 8'b1110001;
DRAM[2899] = 8'b1110001;
DRAM[2900] = 8'b1110010;
DRAM[2901] = 8'b1110010;
DRAM[2902] = 8'b1110010;
DRAM[2903] = 8'b1110010;
DRAM[2904] = 8'b1110000;
DRAM[2905] = 8'b1110000;
DRAM[2906] = 8'b1110000;
DRAM[2907] = 8'b1110000;
DRAM[2908] = 8'b1110000;
DRAM[2909] = 8'b1110000;
DRAM[2910] = 8'b1110000;
DRAM[2911] = 8'b1110000;
DRAM[2912] = 8'b1110010;
DRAM[2913] = 8'b1110001;
DRAM[2914] = 8'b1101111;
DRAM[2915] = 8'b1110000;
DRAM[2916] = 8'b1110010;
DRAM[2917] = 8'b1110010;
DRAM[2918] = 8'b1110001;
DRAM[2919] = 8'b1110000;
DRAM[2920] = 8'b1101111;
DRAM[2921] = 8'b1101111;
DRAM[2922] = 8'b1110000;
DRAM[2923] = 8'b1110000;
DRAM[2924] = 8'b1110000;
DRAM[2925] = 8'b1110000;
DRAM[2926] = 8'b1101111;
DRAM[2927] = 8'b1101111;
DRAM[2928] = 8'b1101111;
DRAM[2929] = 8'b1101111;
DRAM[2930] = 8'b1101111;
DRAM[2931] = 8'b1101111;
DRAM[2932] = 8'b1101111;
DRAM[2933] = 8'b1101111;
DRAM[2934] = 8'b1101111;
DRAM[2935] = 8'b1101111;
DRAM[2936] = 8'b1101111;
DRAM[2937] = 8'b1101111;
DRAM[2938] = 8'b1101111;
DRAM[2939] = 8'b1101111;
DRAM[2940] = 8'b1101111;
DRAM[2941] = 8'b1101111;
DRAM[2942] = 8'b1101111;
DRAM[2943] = 8'b1101111;
DRAM[2944] = 8'b1101111;
DRAM[2945] = 8'b1101111;
DRAM[2946] = 8'b1101111;
DRAM[2947] = 8'b1101111;
DRAM[2948] = 8'b1101111;
DRAM[2949] = 8'b1101111;
DRAM[2950] = 8'b1101111;
DRAM[2951] = 8'b1101111;
DRAM[2952] = 8'b1101111;
DRAM[2953] = 8'b1110000;
DRAM[2954] = 8'b1110001;
DRAM[2955] = 8'b1110001;
DRAM[2956] = 8'b1110001;
DRAM[2957] = 8'b1110001;
DRAM[2958] = 8'b1110000;
DRAM[2959] = 8'b1101111;
DRAM[2960] = 8'b1101110;
DRAM[2961] = 8'b1101110;
DRAM[2962] = 8'b1101111;
DRAM[2963] = 8'b1101111;
DRAM[2964] = 8'b1101111;
DRAM[2965] = 8'b1101111;
DRAM[2966] = 8'b1101110;
DRAM[2967] = 8'b1101110;
DRAM[2968] = 8'b1101110;
DRAM[2969] = 8'b1101110;
DRAM[2970] = 8'b1101110;
DRAM[2971] = 8'b1101110;
DRAM[2972] = 8'b1101110;
DRAM[2973] = 8'b1101110;
DRAM[2974] = 8'b1101110;
DRAM[2975] = 8'b1101110;
DRAM[2976] = 8'b1101100;
DRAM[2977] = 8'b1101100;
DRAM[2978] = 8'b1101100;
DRAM[2979] = 8'b1101100;
DRAM[2980] = 8'b1101011;
DRAM[2981] = 8'b1101011;
DRAM[2982] = 8'b1101011;
DRAM[2983] = 8'b1101011;
DRAM[2984] = 8'b1101011;
DRAM[2985] = 8'b1101011;
DRAM[2986] = 8'b1101010;
DRAM[2987] = 8'b1101010;
DRAM[2988] = 8'b1101010;
DRAM[2989] = 8'b1101001;
DRAM[2990] = 8'b1101001;
DRAM[2991] = 8'b1101001;
DRAM[2992] = 8'b1101000;
DRAM[2993] = 8'b1100111;
DRAM[2994] = 8'b1100111;
DRAM[2995] = 8'b1100110;
DRAM[2996] = 8'b1100101;
DRAM[2997] = 8'b1100100;
DRAM[2998] = 8'b1100100;
DRAM[2999] = 8'b1100100;
DRAM[3000] = 8'b1100011;
DRAM[3001] = 8'b1100010;
DRAM[3002] = 8'b1100010;
DRAM[3003] = 8'b1100001;
DRAM[3004] = 8'b1100000;
DRAM[3005] = 8'b1011111;
DRAM[3006] = 8'b1011111;
DRAM[3007] = 8'b1011111;
DRAM[3008] = 8'b1011110;
DRAM[3009] = 8'b1011101;
DRAM[3010] = 8'b1011101;
DRAM[3011] = 8'b1011100;
DRAM[3012] = 8'b1011011;
DRAM[3013] = 8'b1011010;
DRAM[3014] = 8'b1011010;
DRAM[3015] = 8'b1011010;
DRAM[3016] = 8'b1011000;
DRAM[3017] = 8'b1011000;
DRAM[3018] = 8'b1011000;
DRAM[3019] = 8'b1011000;
DRAM[3020] = 8'b1011000;
DRAM[3021] = 8'b1011000;
DRAM[3022] = 8'b1010111;
DRAM[3023] = 8'b1010111;
DRAM[3024] = 8'b1010110;
DRAM[3025] = 8'b1010101;
DRAM[3026] = 8'b1010100;
DRAM[3027] = 8'b1010010;
DRAM[3028] = 8'b1010010;
DRAM[3029] = 8'b1010001;
DRAM[3030] = 8'b1010001;
DRAM[3031] = 8'b1010010;
DRAM[3032] = 8'b1001111;
DRAM[3033] = 8'b1001111;
DRAM[3034] = 8'b1001111;
DRAM[3035] = 8'b1001111;
DRAM[3036] = 8'b1001111;
DRAM[3037] = 8'b1001111;
DRAM[3038] = 8'b1001111;
DRAM[3039] = 8'b1001111;
DRAM[3040] = 8'b1001110;
DRAM[3041] = 8'b1001101;
DRAM[3042] = 8'b1001100;
DRAM[3043] = 8'b1001011;
DRAM[3044] = 8'b1001011;
DRAM[3045] = 8'b1001011;
DRAM[3046] = 8'b1001011;
DRAM[3047] = 8'b1001100;
DRAM[3048] = 8'b1001010;
DRAM[3049] = 8'b1001010;
DRAM[3050] = 8'b1001001;
DRAM[3051] = 8'b1001001;
DRAM[3052] = 8'b1001000;
DRAM[3053] = 8'b1001000;
DRAM[3054] = 8'b1000111;
DRAM[3055] = 8'b1000111;
DRAM[3056] = 8'b1000111;
DRAM[3057] = 8'b1000110;
DRAM[3058] = 8'b1000110;
DRAM[3059] = 8'b1000110;
DRAM[3060] = 8'b1000101;
DRAM[3061] = 8'b1000101;
DRAM[3062] = 8'b1000101;
DRAM[3063] = 8'b1000101;
DRAM[3064] = 8'b1000011;
DRAM[3065] = 8'b1000011;
DRAM[3066] = 8'b1000010;
DRAM[3067] = 8'b1000010;
DRAM[3068] = 8'b1000010;
DRAM[3069] = 8'b1000001;
DRAM[3070] = 8'b1000001;
DRAM[3071] = 8'b1000001;
DRAM[3072] = 8'b1011111;
DRAM[3073] = 8'b1011111;
DRAM[3074] = 8'b1011111;
DRAM[3075] = 8'b1100000;
DRAM[3076] = 8'b1100001;
DRAM[3077] = 8'b1100001;
DRAM[3078] = 8'b1100010;
DRAM[3079] = 8'b1100010;
DRAM[3080] = 8'b1100011;
DRAM[3081] = 8'b1100011;
DRAM[3082] = 8'b1100011;
DRAM[3083] = 8'b1100011;
DRAM[3084] = 8'b1100011;
DRAM[3085] = 8'b1100100;
DRAM[3086] = 8'b1100100;
DRAM[3087] = 8'b1100100;
DRAM[3088] = 8'b1100101;
DRAM[3089] = 8'b1100101;
DRAM[3090] = 8'b1100110;
DRAM[3091] = 8'b1100110;
DRAM[3092] = 8'b1100111;
DRAM[3093] = 8'b1101000;
DRAM[3094] = 8'b1101001;
DRAM[3095] = 8'b1101001;
DRAM[3096] = 8'b1100110;
DRAM[3097] = 8'b1100111;
DRAM[3098] = 8'b1101000;
DRAM[3099] = 8'b1101001;
DRAM[3100] = 8'b1101001;
DRAM[3101] = 8'b1101001;
DRAM[3102] = 8'b1101001;
DRAM[3103] = 8'b1101001;
DRAM[3104] = 8'b1101011;
DRAM[3105] = 8'b1101100;
DRAM[3106] = 8'b1101100;
DRAM[3107] = 8'b1101100;
DRAM[3108] = 8'b1101101;
DRAM[3109] = 8'b1101101;
DRAM[3110] = 8'b1101101;
DRAM[3111] = 8'b1101110;
DRAM[3112] = 8'b1101101;
DRAM[3113] = 8'b1101101;
DRAM[3114] = 8'b1101110;
DRAM[3115] = 8'b1101110;
DRAM[3116] = 8'b1101110;
DRAM[3117] = 8'b1101111;
DRAM[3118] = 8'b1101111;
DRAM[3119] = 8'b1101111;
DRAM[3120] = 8'b1110001;
DRAM[3121] = 8'b1110001;
DRAM[3122] = 8'b1110010;
DRAM[3123] = 8'b1110010;
DRAM[3124] = 8'b1110011;
DRAM[3125] = 8'b1110011;
DRAM[3126] = 8'b1110011;
DRAM[3127] = 8'b1110011;
DRAM[3128] = 8'b1110100;
DRAM[3129] = 8'b1110100;
DRAM[3130] = 8'b1110100;
DRAM[3131] = 8'b1110100;
DRAM[3132] = 8'b1110100;
DRAM[3133] = 8'b1110100;
DRAM[3134] = 8'b1110100;
DRAM[3135] = 8'b1110100;
DRAM[3136] = 8'b1110011;
DRAM[3137] = 8'b1110011;
DRAM[3138] = 8'b1110011;
DRAM[3139] = 8'b1110011;
DRAM[3140] = 8'b1110011;
DRAM[3141] = 8'b1110011;
DRAM[3142] = 8'b1110011;
DRAM[3143] = 8'b1110011;
DRAM[3144] = 8'b1110010;
DRAM[3145] = 8'b1110010;
DRAM[3146] = 8'b1110010;
DRAM[3147] = 8'b1110010;
DRAM[3148] = 8'b1110010;
DRAM[3149] = 8'b1110010;
DRAM[3150] = 8'b1110010;
DRAM[3151] = 8'b1110010;
DRAM[3152] = 8'b1110010;
DRAM[3153] = 8'b1110010;
DRAM[3154] = 8'b1110010;
DRAM[3155] = 8'b1110010;
DRAM[3156] = 8'b1110011;
DRAM[3157] = 8'b1110011;
DRAM[3158] = 8'b1110011;
DRAM[3159] = 8'b1110011;
DRAM[3160] = 8'b1110000;
DRAM[3161] = 8'b1110000;
DRAM[3162] = 8'b1110000;
DRAM[3163] = 8'b1110000;
DRAM[3164] = 8'b1110000;
DRAM[3165] = 8'b1110000;
DRAM[3166] = 8'b1110000;
DRAM[3167] = 8'b1110000;
DRAM[3168] = 8'b1110010;
DRAM[3169] = 8'b1110001;
DRAM[3170] = 8'b1110000;
DRAM[3171] = 8'b1110000;
DRAM[3172] = 8'b1110010;
DRAM[3173] = 8'b1110011;
DRAM[3174] = 8'b1110001;
DRAM[3175] = 8'b1110000;
DRAM[3176] = 8'b1101111;
DRAM[3177] = 8'b1110000;
DRAM[3178] = 8'b1110000;
DRAM[3179] = 8'b1110001;
DRAM[3180] = 8'b1110001;
DRAM[3181] = 8'b1110000;
DRAM[3182] = 8'b1110000;
DRAM[3183] = 8'b1101111;
DRAM[3184] = 8'b1101111;
DRAM[3185] = 8'b1101111;
DRAM[3186] = 8'b1101111;
DRAM[3187] = 8'b1101111;
DRAM[3188] = 8'b1101111;
DRAM[3189] = 8'b1101111;
DRAM[3190] = 8'b1101111;
DRAM[3191] = 8'b1101111;
DRAM[3192] = 8'b1101111;
DRAM[3193] = 8'b1101111;
DRAM[3194] = 8'b1101111;
DRAM[3195] = 8'b1101111;
DRAM[3196] = 8'b1101111;
DRAM[3197] = 8'b1101111;
DRAM[3198] = 8'b1101111;
DRAM[3199] = 8'b1101111;
DRAM[3200] = 8'b1101111;
DRAM[3201] = 8'b1101111;
DRAM[3202] = 8'b1101111;
DRAM[3203] = 8'b1101111;
DRAM[3204] = 8'b1101111;
DRAM[3205] = 8'b1101111;
DRAM[3206] = 8'b1101111;
DRAM[3207] = 8'b1101111;
DRAM[3208] = 8'b1101111;
DRAM[3209] = 8'b1101111;
DRAM[3210] = 8'b1110000;
DRAM[3211] = 8'b1110001;
DRAM[3212] = 8'b1110001;
DRAM[3213] = 8'b1110000;
DRAM[3214] = 8'b1101111;
DRAM[3215] = 8'b1101111;
DRAM[3216] = 8'b1101110;
DRAM[3217] = 8'b1101111;
DRAM[3218] = 8'b1110000;
DRAM[3219] = 8'b1110000;
DRAM[3220] = 8'b1110000;
DRAM[3221] = 8'b1110000;
DRAM[3222] = 8'b1101111;
DRAM[3223] = 8'b1101110;
DRAM[3224] = 8'b1101110;
DRAM[3225] = 8'b1101110;
DRAM[3226] = 8'b1101110;
DRAM[3227] = 8'b1101110;
DRAM[3228] = 8'b1101110;
DRAM[3229] = 8'b1101110;
DRAM[3230] = 8'b1101110;
DRAM[3231] = 8'b1101110;
DRAM[3232] = 8'b1101110;
DRAM[3233] = 8'b1101110;
DRAM[3234] = 8'b1101101;
DRAM[3235] = 8'b1101101;
DRAM[3236] = 8'b1101100;
DRAM[3237] = 8'b1101100;
DRAM[3238] = 8'b1101011;
DRAM[3239] = 8'b1101011;
DRAM[3240] = 8'b1101100;
DRAM[3241] = 8'b1101011;
DRAM[3242] = 8'b1101011;
DRAM[3243] = 8'b1101011;
DRAM[3244] = 8'b1101010;
DRAM[3245] = 8'b1101010;
DRAM[3246] = 8'b1101010;
DRAM[3247] = 8'b1101010;
DRAM[3248] = 8'b1101000;
DRAM[3249] = 8'b1101000;
DRAM[3250] = 8'b1101000;
DRAM[3251] = 8'b1100111;
DRAM[3252] = 8'b1100110;
DRAM[3253] = 8'b1100101;
DRAM[3254] = 8'b1100101;
DRAM[3255] = 8'b1100100;
DRAM[3256] = 8'b1100011;
DRAM[3257] = 8'b1100011;
DRAM[3258] = 8'b1100011;
DRAM[3259] = 8'b1100010;
DRAM[3260] = 8'b1100001;
DRAM[3261] = 8'b1100000;
DRAM[3262] = 8'b1100000;
DRAM[3263] = 8'b1011111;
DRAM[3264] = 8'b1011110;
DRAM[3265] = 8'b1011110;
DRAM[3266] = 8'b1011110;
DRAM[3267] = 8'b1011101;
DRAM[3268] = 8'b1011100;
DRAM[3269] = 8'b1011011;
DRAM[3270] = 8'b1011011;
DRAM[3271] = 8'b1011010;
DRAM[3272] = 8'b1011001;
DRAM[3273] = 8'b1011001;
DRAM[3274] = 8'b1011000;
DRAM[3275] = 8'b1011000;
DRAM[3276] = 8'b1011000;
DRAM[3277] = 8'b1011000;
DRAM[3278] = 8'b1011000;
DRAM[3279] = 8'b1011000;
DRAM[3280] = 8'b1010110;
DRAM[3281] = 8'b1010101;
DRAM[3282] = 8'b1010100;
DRAM[3283] = 8'b1010011;
DRAM[3284] = 8'b1010010;
DRAM[3285] = 8'b1010010;
DRAM[3286] = 8'b1010010;
DRAM[3287] = 8'b1010010;
DRAM[3288] = 8'b1001111;
DRAM[3289] = 8'b1001111;
DRAM[3290] = 8'b1001111;
DRAM[3291] = 8'b1001111;
DRAM[3292] = 8'b1001111;
DRAM[3293] = 8'b1001111;
DRAM[3294] = 8'b1001111;
DRAM[3295] = 8'b1001111;
DRAM[3296] = 8'b1001110;
DRAM[3297] = 8'b1001101;
DRAM[3298] = 8'b1001100;
DRAM[3299] = 8'b1001100;
DRAM[3300] = 8'b1001011;
DRAM[3301] = 8'b1001011;
DRAM[3302] = 8'b1001100;
DRAM[3303] = 8'b1001100;
DRAM[3304] = 8'b1001010;
DRAM[3305] = 8'b1001010;
DRAM[3306] = 8'b1001010;
DRAM[3307] = 8'b1001010;
DRAM[3308] = 8'b1001001;
DRAM[3309] = 8'b1001001;
DRAM[3310] = 8'b1001001;
DRAM[3311] = 8'b1001001;
DRAM[3312] = 8'b1000111;
DRAM[3313] = 8'b1000111;
DRAM[3314] = 8'b1000111;
DRAM[3315] = 8'b1000111;
DRAM[3316] = 8'b1000110;
DRAM[3317] = 8'b1000110;
DRAM[3318] = 8'b1000110;
DRAM[3319] = 8'b1000101;
DRAM[3320] = 8'b1000011;
DRAM[3321] = 8'b1000011;
DRAM[3322] = 8'b1000011;
DRAM[3323] = 8'b1000010;
DRAM[3324] = 8'b1000010;
DRAM[3325] = 8'b1000010;
DRAM[3326] = 8'b1000001;
DRAM[3327] = 8'b1000001;
DRAM[3328] = 8'b1100000;
DRAM[3329] = 8'b1100000;
DRAM[3330] = 8'b1100000;
DRAM[3331] = 8'b1100001;
DRAM[3332] = 8'b1100001;
DRAM[3333] = 8'b1100010;
DRAM[3334] = 8'b1100010;
DRAM[3335] = 8'b1100010;
DRAM[3336] = 8'b1100011;
DRAM[3337] = 8'b1100011;
DRAM[3338] = 8'b1100011;
DRAM[3339] = 8'b1100011;
DRAM[3340] = 8'b1100011;
DRAM[3341] = 8'b1100011;
DRAM[3342] = 8'b1100011;
DRAM[3343] = 8'b1100011;
DRAM[3344] = 8'b1100110;
DRAM[3345] = 8'b1100110;
DRAM[3346] = 8'b1100111;
DRAM[3347] = 8'b1100111;
DRAM[3348] = 8'b1101000;
DRAM[3349] = 8'b1101001;
DRAM[3350] = 8'b1101010;
DRAM[3351] = 8'b1101010;
DRAM[3352] = 8'b1101000;
DRAM[3353] = 8'b1101000;
DRAM[3354] = 8'b1101001;
DRAM[3355] = 8'b1101010;
DRAM[3356] = 8'b1101011;
DRAM[3357] = 8'b1101011;
DRAM[3358] = 8'b1101010;
DRAM[3359] = 8'b1101010;
DRAM[3360] = 8'b1101011;
DRAM[3361] = 8'b1101011;
DRAM[3362] = 8'b1101100;
DRAM[3363] = 8'b1101100;
DRAM[3364] = 8'b1101101;
DRAM[3365] = 8'b1101101;
DRAM[3366] = 8'b1101101;
DRAM[3367] = 8'b1101101;
DRAM[3368] = 8'b1101110;
DRAM[3369] = 8'b1101110;
DRAM[3370] = 8'b1101110;
DRAM[3371] = 8'b1101110;
DRAM[3372] = 8'b1101111;
DRAM[3373] = 8'b1101111;
DRAM[3374] = 8'b1101111;
DRAM[3375] = 8'b1110000;
DRAM[3376] = 8'b1110001;
DRAM[3377] = 8'b1110001;
DRAM[3378] = 8'b1110010;
DRAM[3379] = 8'b1110011;
DRAM[3380] = 8'b1110100;
DRAM[3381] = 8'b1110100;
DRAM[3382] = 8'b1110011;
DRAM[3383] = 8'b1110011;
DRAM[3384] = 8'b1110100;
DRAM[3385] = 8'b1110100;
DRAM[3386] = 8'b1110100;
DRAM[3387] = 8'b1110100;
DRAM[3388] = 8'b1110100;
DRAM[3389] = 8'b1110100;
DRAM[3390] = 8'b1110100;
DRAM[3391] = 8'b1110100;
DRAM[3392] = 8'b1110100;
DRAM[3393] = 8'b1110100;
DRAM[3394] = 8'b1110100;
DRAM[3395] = 8'b1110100;
DRAM[3396] = 8'b1110100;
DRAM[3397] = 8'b1110100;
DRAM[3398] = 8'b1110100;
DRAM[3399] = 8'b1110100;
DRAM[3400] = 8'b1110011;
DRAM[3401] = 8'b1110011;
DRAM[3402] = 8'b1110011;
DRAM[3403] = 8'b1110011;
DRAM[3404] = 8'b1110011;
DRAM[3405] = 8'b1110011;
DRAM[3406] = 8'b1110011;
DRAM[3407] = 8'b1110011;
DRAM[3408] = 8'b1110100;
DRAM[3409] = 8'b1110100;
DRAM[3410] = 8'b1110011;
DRAM[3411] = 8'b1110011;
DRAM[3412] = 8'b1110011;
DRAM[3413] = 8'b1110011;
DRAM[3414] = 8'b1110011;
DRAM[3415] = 8'b1110011;
DRAM[3416] = 8'b1110001;
DRAM[3417] = 8'b1110001;
DRAM[3418] = 8'b1110001;
DRAM[3419] = 8'b1110001;
DRAM[3420] = 8'b1110001;
DRAM[3421] = 8'b1110001;
DRAM[3422] = 8'b1110001;
DRAM[3423] = 8'b1110001;
DRAM[3424] = 8'b1110011;
DRAM[3425] = 8'b1110001;
DRAM[3426] = 8'b1110000;
DRAM[3427] = 8'b1110001;
DRAM[3428] = 8'b1110010;
DRAM[3429] = 8'b1110011;
DRAM[3430] = 8'b1110010;
DRAM[3431] = 8'b1110000;
DRAM[3432] = 8'b1110000;
DRAM[3433] = 8'b1110001;
DRAM[3434] = 8'b1110001;
DRAM[3435] = 8'b1110010;
DRAM[3436] = 8'b1110010;
DRAM[3437] = 8'b1110001;
DRAM[3438] = 8'b1110001;
DRAM[3439] = 8'b1110000;
DRAM[3440] = 8'b1110000;
DRAM[3441] = 8'b1110000;
DRAM[3442] = 8'b1110000;
DRAM[3443] = 8'b1110000;
DRAM[3444] = 8'b1110000;
DRAM[3445] = 8'b1110000;
DRAM[3446] = 8'b1110000;
DRAM[3447] = 8'b1110000;
DRAM[3448] = 8'b1110000;
DRAM[3449] = 8'b1110000;
DRAM[3450] = 8'b1110000;
DRAM[3451] = 8'b1110000;
DRAM[3452] = 8'b1110000;
DRAM[3453] = 8'b1110000;
DRAM[3454] = 8'b1110000;
DRAM[3455] = 8'b1110000;
DRAM[3456] = 8'b1110000;
DRAM[3457] = 8'b1110000;
DRAM[3458] = 8'b1110000;
DRAM[3459] = 8'b1110000;
DRAM[3460] = 8'b1110000;
DRAM[3461] = 8'b1110000;
DRAM[3462] = 8'b1110000;
DRAM[3463] = 8'b1110000;
DRAM[3464] = 8'b1101111;
DRAM[3465] = 8'b1110000;
DRAM[3466] = 8'b1110000;
DRAM[3467] = 8'b1110001;
DRAM[3468] = 8'b1110001;
DRAM[3469] = 8'b1110000;
DRAM[3470] = 8'b1110000;
DRAM[3471] = 8'b1101111;
DRAM[3472] = 8'b1110000;
DRAM[3473] = 8'b1110000;
DRAM[3474] = 8'b1110001;
DRAM[3475] = 8'b1110010;
DRAM[3476] = 8'b1110010;
DRAM[3477] = 8'b1110001;
DRAM[3478] = 8'b1110000;
DRAM[3479] = 8'b1110000;
DRAM[3480] = 8'b1101111;
DRAM[3481] = 8'b1101111;
DRAM[3482] = 8'b1101111;
DRAM[3483] = 8'b1101111;
DRAM[3484] = 8'b1101111;
DRAM[3485] = 8'b1101111;
DRAM[3486] = 8'b1101111;
DRAM[3487] = 8'b1101111;
DRAM[3488] = 8'b1101111;
DRAM[3489] = 8'b1101111;
DRAM[3490] = 8'b1101110;
DRAM[3491] = 8'b1101110;
DRAM[3492] = 8'b1101101;
DRAM[3493] = 8'b1101100;
DRAM[3494] = 8'b1101100;
DRAM[3495] = 8'b1101011;
DRAM[3496] = 8'b1101100;
DRAM[3497] = 8'b1101100;
DRAM[3498] = 8'b1101011;
DRAM[3499] = 8'b1101011;
DRAM[3500] = 8'b1101010;
DRAM[3501] = 8'b1101010;
DRAM[3502] = 8'b1101010;
DRAM[3503] = 8'b1101010;
DRAM[3504] = 8'b1101001;
DRAM[3505] = 8'b1101001;
DRAM[3506] = 8'b1101000;
DRAM[3507] = 8'b1101000;
DRAM[3508] = 8'b1100111;
DRAM[3509] = 8'b1100110;
DRAM[3510] = 8'b1100101;
DRAM[3511] = 8'b1100101;
DRAM[3512] = 8'b1100100;
DRAM[3513] = 8'b1100100;
DRAM[3514] = 8'b1100011;
DRAM[3515] = 8'b1100011;
DRAM[3516] = 8'b1100010;
DRAM[3517] = 8'b1100001;
DRAM[3518] = 8'b1100000;
DRAM[3519] = 8'b1100000;
DRAM[3520] = 8'b1011111;
DRAM[3521] = 8'b1011111;
DRAM[3522] = 8'b1011110;
DRAM[3523] = 8'b1011110;
DRAM[3524] = 8'b1011101;
DRAM[3525] = 8'b1011100;
DRAM[3526] = 8'b1011011;
DRAM[3527] = 8'b1011011;
DRAM[3528] = 8'b1011010;
DRAM[3529] = 8'b1011010;
DRAM[3530] = 8'b1011001;
DRAM[3531] = 8'b1011001;
DRAM[3532] = 8'b1011000;
DRAM[3533] = 8'b1011000;
DRAM[3534] = 8'b1010111;
DRAM[3535] = 8'b1010111;
DRAM[3536] = 8'b1010110;
DRAM[3537] = 8'b1010110;
DRAM[3538] = 8'b1010100;
DRAM[3539] = 8'b1010011;
DRAM[3540] = 8'b1010010;
DRAM[3541] = 8'b1010010;
DRAM[3542] = 8'b1010010;
DRAM[3543] = 8'b1010010;
DRAM[3544] = 8'b1001111;
DRAM[3545] = 8'b1001111;
DRAM[3546] = 8'b1001111;
DRAM[3547] = 8'b1001111;
DRAM[3548] = 8'b1001111;
DRAM[3549] = 8'b1001111;
DRAM[3550] = 8'b1001111;
DRAM[3551] = 8'b1001111;
DRAM[3552] = 8'b1001110;
DRAM[3553] = 8'b1001110;
DRAM[3554] = 8'b1001101;
DRAM[3555] = 8'b1001100;
DRAM[3556] = 8'b1001100;
DRAM[3557] = 8'b1001100;
DRAM[3558] = 8'b1001100;
DRAM[3559] = 8'b1001100;
DRAM[3560] = 8'b1001010;
DRAM[3561] = 8'b1001010;
DRAM[3562] = 8'b1001010;
DRAM[3563] = 8'b1001010;
DRAM[3564] = 8'b1001010;
DRAM[3565] = 8'b1001010;
DRAM[3566] = 8'b1001010;
DRAM[3567] = 8'b1001010;
DRAM[3568] = 8'b1001000;
DRAM[3569] = 8'b1001000;
DRAM[3570] = 8'b1001000;
DRAM[3571] = 8'b1000111;
DRAM[3572] = 8'b1000111;
DRAM[3573] = 8'b1000111;
DRAM[3574] = 8'b1000110;
DRAM[3575] = 8'b1000110;
DRAM[3576] = 8'b1000100;
DRAM[3577] = 8'b1000011;
DRAM[3578] = 8'b1000011;
DRAM[3579] = 8'b1000011;
DRAM[3580] = 8'b1000010;
DRAM[3581] = 8'b1000010;
DRAM[3582] = 8'b1000010;
DRAM[3583] = 8'b1000010;
DRAM[3584] = 8'b1100001;
DRAM[3585] = 8'b1100001;
DRAM[3586] = 8'b1100001;
DRAM[3587] = 8'b1100010;
DRAM[3588] = 8'b1100010;
DRAM[3589] = 8'b1100010;
DRAM[3590] = 8'b1100010;
DRAM[3591] = 8'b1100011;
DRAM[3592] = 8'b1100100;
DRAM[3593] = 8'b1100100;
DRAM[3594] = 8'b1100100;
DRAM[3595] = 8'b1100100;
DRAM[3596] = 8'b1100100;
DRAM[3597] = 8'b1100100;
DRAM[3598] = 8'b1100100;
DRAM[3599] = 8'b1100100;
DRAM[3600] = 8'b1100101;
DRAM[3601] = 8'b1100101;
DRAM[3602] = 8'b1100110;
DRAM[3603] = 8'b1100111;
DRAM[3604] = 8'b1101000;
DRAM[3605] = 8'b1101000;
DRAM[3606] = 8'b1101001;
DRAM[3607] = 8'b1101001;
DRAM[3608] = 8'b1101001;
DRAM[3609] = 8'b1101010;
DRAM[3610] = 8'b1101011;
DRAM[3611] = 8'b1101100;
DRAM[3612] = 8'b1101100;
DRAM[3613] = 8'b1101100;
DRAM[3614] = 8'b1101100;
DRAM[3615] = 8'b1101011;
DRAM[3616] = 8'b1101101;
DRAM[3617] = 8'b1101101;
DRAM[3618] = 8'b1101101;
DRAM[3619] = 8'b1101101;
DRAM[3620] = 8'b1101110;
DRAM[3621] = 8'b1101110;
DRAM[3622] = 8'b1101111;
DRAM[3623] = 8'b1101111;
DRAM[3624] = 8'b1101110;
DRAM[3625] = 8'b1101110;
DRAM[3626] = 8'b1101110;
DRAM[3627] = 8'b1101111;
DRAM[3628] = 8'b1101111;
DRAM[3629] = 8'b1101111;
DRAM[3630] = 8'b1110000;
DRAM[3631] = 8'b1110000;
DRAM[3632] = 8'b1110000;
DRAM[3633] = 8'b1110001;
DRAM[3634] = 8'b1110011;
DRAM[3635] = 8'b1110100;
DRAM[3636] = 8'b1110100;
DRAM[3637] = 8'b1110100;
DRAM[3638] = 8'b1110011;
DRAM[3639] = 8'b1110011;
DRAM[3640] = 8'b1110011;
DRAM[3641] = 8'b1110011;
DRAM[3642] = 8'b1110011;
DRAM[3643] = 8'b1110011;
DRAM[3644] = 8'b1110011;
DRAM[3645] = 8'b1110011;
DRAM[3646] = 8'b1110011;
DRAM[3647] = 8'b1110011;
DRAM[3648] = 8'b1110100;
DRAM[3649] = 8'b1110100;
DRAM[3650] = 8'b1110100;
DRAM[3651] = 8'b1110100;
DRAM[3652] = 8'b1110100;
DRAM[3653] = 8'b1110100;
DRAM[3654] = 8'b1110100;
DRAM[3655] = 8'b1110100;
DRAM[3656] = 8'b1110011;
DRAM[3657] = 8'b1110011;
DRAM[3658] = 8'b1110011;
DRAM[3659] = 8'b1110011;
DRAM[3660] = 8'b1110011;
DRAM[3661] = 8'b1110011;
DRAM[3662] = 8'b1110011;
DRAM[3663] = 8'b1110011;
DRAM[3664] = 8'b1110101;
DRAM[3665] = 8'b1110101;
DRAM[3666] = 8'b1110101;
DRAM[3667] = 8'b1110100;
DRAM[3668] = 8'b1110011;
DRAM[3669] = 8'b1110011;
DRAM[3670] = 8'b1110010;
DRAM[3671] = 8'b1110010;
DRAM[3672] = 8'b1110001;
DRAM[3673] = 8'b1110001;
DRAM[3674] = 8'b1110001;
DRAM[3675] = 8'b1110001;
DRAM[3676] = 8'b1110001;
DRAM[3677] = 8'b1110001;
DRAM[3678] = 8'b1110001;
DRAM[3679] = 8'b1110001;
DRAM[3680] = 8'b1110011;
DRAM[3681] = 8'b1110010;
DRAM[3682] = 8'b1110000;
DRAM[3683] = 8'b1110001;
DRAM[3684] = 8'b1110011;
DRAM[3685] = 8'b1110011;
DRAM[3686] = 8'b1110010;
DRAM[3687] = 8'b1110001;
DRAM[3688] = 8'b1110010;
DRAM[3689] = 8'b1110010;
DRAM[3690] = 8'b1110011;
DRAM[3691] = 8'b1110011;
DRAM[3692] = 8'b1110011;
DRAM[3693] = 8'b1110011;
DRAM[3694] = 8'b1110010;
DRAM[3695] = 8'b1110010;
DRAM[3696] = 8'b1110001;
DRAM[3697] = 8'b1110001;
DRAM[3698] = 8'b1110001;
DRAM[3699] = 8'b1110001;
DRAM[3700] = 8'b1110001;
DRAM[3701] = 8'b1110001;
DRAM[3702] = 8'b1110001;
DRAM[3703] = 8'b1110001;
DRAM[3704] = 8'b1110001;
DRAM[3705] = 8'b1110001;
DRAM[3706] = 8'b1110001;
DRAM[3707] = 8'b1110001;
DRAM[3708] = 8'b1110001;
DRAM[3709] = 8'b1110001;
DRAM[3710] = 8'b1110001;
DRAM[3711] = 8'b1110001;
DRAM[3712] = 8'b1110001;
DRAM[3713] = 8'b1110001;
DRAM[3714] = 8'b1110001;
DRAM[3715] = 8'b1110001;
DRAM[3716] = 8'b1110001;
DRAM[3717] = 8'b1110001;
DRAM[3718] = 8'b1110001;
DRAM[3719] = 8'b1110001;
DRAM[3720] = 8'b1110001;
DRAM[3721] = 8'b1110001;
DRAM[3722] = 8'b1110010;
DRAM[3723] = 8'b1110010;
DRAM[3724] = 8'b1110010;
DRAM[3725] = 8'b1110010;
DRAM[3726] = 8'b1110001;
DRAM[3727] = 8'b1110001;
DRAM[3728] = 8'b1110001;
DRAM[3729] = 8'b1110010;
DRAM[3730] = 8'b1110011;
DRAM[3731] = 8'b1110011;
DRAM[3732] = 8'b1110011;
DRAM[3733] = 8'b1110011;
DRAM[3734] = 8'b1110010;
DRAM[3735] = 8'b1110001;
DRAM[3736] = 8'b1110000;
DRAM[3737] = 8'b1110000;
DRAM[3738] = 8'b1110000;
DRAM[3739] = 8'b1110000;
DRAM[3740] = 8'b1110000;
DRAM[3741] = 8'b1110000;
DRAM[3742] = 8'b1110000;
DRAM[3743] = 8'b1110000;
DRAM[3744] = 8'b1110000;
DRAM[3745] = 8'b1110000;
DRAM[3746] = 8'b1101111;
DRAM[3747] = 8'b1101110;
DRAM[3748] = 8'b1101101;
DRAM[3749] = 8'b1101100;
DRAM[3750] = 8'b1101100;
DRAM[3751] = 8'b1101011;
DRAM[3752] = 8'b1101011;
DRAM[3753] = 8'b1101011;
DRAM[3754] = 8'b1101011;
DRAM[3755] = 8'b1101010;
DRAM[3756] = 8'b1101010;
DRAM[3757] = 8'b1101010;
DRAM[3758] = 8'b1101001;
DRAM[3759] = 8'b1101001;
DRAM[3760] = 8'b1101010;
DRAM[3761] = 8'b1101010;
DRAM[3762] = 8'b1101001;
DRAM[3763] = 8'b1101000;
DRAM[3764] = 8'b1100111;
DRAM[3765] = 8'b1100111;
DRAM[3766] = 8'b1100110;
DRAM[3767] = 8'b1100110;
DRAM[3768] = 8'b1100101;
DRAM[3769] = 8'b1100101;
DRAM[3770] = 8'b1100100;
DRAM[3771] = 8'b1100011;
DRAM[3772] = 8'b1100010;
DRAM[3773] = 8'b1100010;
DRAM[3774] = 8'b1100001;
DRAM[3775] = 8'b1100001;
DRAM[3776] = 8'b1100000;
DRAM[3777] = 8'b1100000;
DRAM[3778] = 8'b1011111;
DRAM[3779] = 8'b1011110;
DRAM[3780] = 8'b1011101;
DRAM[3781] = 8'b1011101;
DRAM[3782] = 8'b1011100;
DRAM[3783] = 8'b1011100;
DRAM[3784] = 8'b1011100;
DRAM[3785] = 8'b1011011;
DRAM[3786] = 8'b1011010;
DRAM[3787] = 8'b1011001;
DRAM[3788] = 8'b1011000;
DRAM[3789] = 8'b1010111;
DRAM[3790] = 8'b1010111;
DRAM[3791] = 8'b1010110;
DRAM[3792] = 8'b1010111;
DRAM[3793] = 8'b1010110;
DRAM[3794] = 8'b1010101;
DRAM[3795] = 8'b1010011;
DRAM[3796] = 8'b1010011;
DRAM[3797] = 8'b1010010;
DRAM[3798] = 8'b1010010;
DRAM[3799] = 8'b1010011;
DRAM[3800] = 8'b1001111;
DRAM[3801] = 8'b1001111;
DRAM[3802] = 8'b1001111;
DRAM[3803] = 8'b1001111;
DRAM[3804] = 8'b1001111;
DRAM[3805] = 8'b1001111;
DRAM[3806] = 8'b1001111;
DRAM[3807] = 8'b1001111;
DRAM[3808] = 8'b1001111;
DRAM[3809] = 8'b1001110;
DRAM[3810] = 8'b1001101;
DRAM[3811] = 8'b1001100;
DRAM[3812] = 8'b1001100;
DRAM[3813] = 8'b1001100;
DRAM[3814] = 8'b1001100;
DRAM[3815] = 8'b1001101;
DRAM[3816] = 8'b1001011;
DRAM[3817] = 8'b1001011;
DRAM[3818] = 8'b1001011;
DRAM[3819] = 8'b1001011;
DRAM[3820] = 8'b1001011;
DRAM[3821] = 8'b1001011;
DRAM[3822] = 8'b1001011;
DRAM[3823] = 8'b1001011;
DRAM[3824] = 8'b1001001;
DRAM[3825] = 8'b1001001;
DRAM[3826] = 8'b1001000;
DRAM[3827] = 8'b1001000;
DRAM[3828] = 8'b1001000;
DRAM[3829] = 8'b1000111;
DRAM[3830] = 8'b1000111;
DRAM[3831] = 8'b1000111;
DRAM[3832] = 8'b1000100;
DRAM[3833] = 8'b1000100;
DRAM[3834] = 8'b1000011;
DRAM[3835] = 8'b1000011;
DRAM[3836] = 8'b1000011;
DRAM[3837] = 8'b1000010;
DRAM[3838] = 8'b1000010;
DRAM[3839] = 8'b1000010;
DRAM[3840] = 8'b1100001;
DRAM[3841] = 8'b1100010;
DRAM[3842] = 8'b1100010;
DRAM[3843] = 8'b1100010;
DRAM[3844] = 8'b1100010;
DRAM[3845] = 8'b1100010;
DRAM[3846] = 8'b1100011;
DRAM[3847] = 8'b1100011;
DRAM[3848] = 8'b1100101;
DRAM[3849] = 8'b1100101;
DRAM[3850] = 8'b1100101;
DRAM[3851] = 8'b1100101;
DRAM[3852] = 8'b1100101;
DRAM[3853] = 8'b1100101;
DRAM[3854] = 8'b1100101;
DRAM[3855] = 8'b1100101;
DRAM[3856] = 8'b1100100;
DRAM[3857] = 8'b1100100;
DRAM[3858] = 8'b1100101;
DRAM[3859] = 8'b1100110;
DRAM[3860] = 8'b1100110;
DRAM[3861] = 8'b1100111;
DRAM[3862] = 8'b1101000;
DRAM[3863] = 8'b1101000;
DRAM[3864] = 8'b1101010;
DRAM[3865] = 8'b1101011;
DRAM[3866] = 8'b1101100;
DRAM[3867] = 8'b1101101;
DRAM[3868] = 8'b1101101;
DRAM[3869] = 8'b1101101;
DRAM[3870] = 8'b1101101;
DRAM[3871] = 8'b1101100;
DRAM[3872] = 8'b1101110;
DRAM[3873] = 8'b1101110;
DRAM[3874] = 8'b1101110;
DRAM[3875] = 8'b1101111;
DRAM[3876] = 8'b1101111;
DRAM[3877] = 8'b1110000;
DRAM[3878] = 8'b1110000;
DRAM[3879] = 8'b1110000;
DRAM[3880] = 8'b1101110;
DRAM[3881] = 8'b1101110;
DRAM[3882] = 8'b1101110;
DRAM[3883] = 8'b1101111;
DRAM[3884] = 8'b1101111;
DRAM[3885] = 8'b1110000;
DRAM[3886] = 8'b1110000;
DRAM[3887] = 8'b1110000;
DRAM[3888] = 8'b1110000;
DRAM[3889] = 8'b1110001;
DRAM[3890] = 8'b1110011;
DRAM[3891] = 8'b1110100;
DRAM[3892] = 8'b1110101;
DRAM[3893] = 8'b1110100;
DRAM[3894] = 8'b1110011;
DRAM[3895] = 8'b1110010;
DRAM[3896] = 8'b1110011;
DRAM[3897] = 8'b1110011;
DRAM[3898] = 8'b1110011;
DRAM[3899] = 8'b1110011;
DRAM[3900] = 8'b1110011;
DRAM[3901] = 8'b1110011;
DRAM[3902] = 8'b1110011;
DRAM[3903] = 8'b1110011;
DRAM[3904] = 8'b1110100;
DRAM[3905] = 8'b1110100;
DRAM[3906] = 8'b1110100;
DRAM[3907] = 8'b1110100;
DRAM[3908] = 8'b1110100;
DRAM[3909] = 8'b1110100;
DRAM[3910] = 8'b1110100;
DRAM[3911] = 8'b1110100;
DRAM[3912] = 8'b1110011;
DRAM[3913] = 8'b1110011;
DRAM[3914] = 8'b1110011;
DRAM[3915] = 8'b1110011;
DRAM[3916] = 8'b1110011;
DRAM[3917] = 8'b1110011;
DRAM[3918] = 8'b1110011;
DRAM[3919] = 8'b1110011;
DRAM[3920] = 8'b1110111;
DRAM[3921] = 8'b1110110;
DRAM[3922] = 8'b1110110;
DRAM[3923] = 8'b1110101;
DRAM[3924] = 8'b1110100;
DRAM[3925] = 8'b1110011;
DRAM[3926] = 8'b1110010;
DRAM[3927] = 8'b1110001;
DRAM[3928] = 8'b1110001;
DRAM[3929] = 8'b1110001;
DRAM[3930] = 8'b1110001;
DRAM[3931] = 8'b1110001;
DRAM[3932] = 8'b1110001;
DRAM[3933] = 8'b1110001;
DRAM[3934] = 8'b1110001;
DRAM[3935] = 8'b1110001;
DRAM[3936] = 8'b1110011;
DRAM[3937] = 8'b1110010;
DRAM[3938] = 8'b1110001;
DRAM[3939] = 8'b1110001;
DRAM[3940] = 8'b1110011;
DRAM[3941] = 8'b1110011;
DRAM[3942] = 8'b1110010;
DRAM[3943] = 8'b1110001;
DRAM[3944] = 8'b1110010;
DRAM[3945] = 8'b1110011;
DRAM[3946] = 8'b1110100;
DRAM[3947] = 8'b1110100;
DRAM[3948] = 8'b1110100;
DRAM[3949] = 8'b1110100;
DRAM[3950] = 8'b1110011;
DRAM[3951] = 8'b1110010;
DRAM[3952] = 8'b1110001;
DRAM[3953] = 8'b1110001;
DRAM[3954] = 8'b1110001;
DRAM[3955] = 8'b1110001;
DRAM[3956] = 8'b1110001;
DRAM[3957] = 8'b1110001;
DRAM[3958] = 8'b1110001;
DRAM[3959] = 8'b1110001;
DRAM[3960] = 8'b1110001;
DRAM[3961] = 8'b1110001;
DRAM[3962] = 8'b1110001;
DRAM[3963] = 8'b1110001;
DRAM[3964] = 8'b1110001;
DRAM[3965] = 8'b1110001;
DRAM[3966] = 8'b1110001;
DRAM[3967] = 8'b1110001;
DRAM[3968] = 8'b1110001;
DRAM[3969] = 8'b1110001;
DRAM[3970] = 8'b1110001;
DRAM[3971] = 8'b1110001;
DRAM[3972] = 8'b1110001;
DRAM[3973] = 8'b1110001;
DRAM[3974] = 8'b1110001;
DRAM[3975] = 8'b1110001;
DRAM[3976] = 8'b1110010;
DRAM[3977] = 8'b1110011;
DRAM[3978] = 8'b1110011;
DRAM[3979] = 8'b1110100;
DRAM[3980] = 8'b1110100;
DRAM[3981] = 8'b1110011;
DRAM[3982] = 8'b1110011;
DRAM[3983] = 8'b1110010;
DRAM[3984] = 8'b1110010;
DRAM[3985] = 8'b1110011;
DRAM[3986] = 8'b1110100;
DRAM[3987] = 8'b1110100;
DRAM[3988] = 8'b1110100;
DRAM[3989] = 8'b1110100;
DRAM[3990] = 8'b1110011;
DRAM[3991] = 8'b1110010;
DRAM[3992] = 8'b1110000;
DRAM[3993] = 8'b1110000;
DRAM[3994] = 8'b1110000;
DRAM[3995] = 8'b1110000;
DRAM[3996] = 8'b1110000;
DRAM[3997] = 8'b1110000;
DRAM[3998] = 8'b1110000;
DRAM[3999] = 8'b1110000;
DRAM[4000] = 8'b1110001;
DRAM[4001] = 8'b1110000;
DRAM[4002] = 8'b1101111;
DRAM[4003] = 8'b1101111;
DRAM[4004] = 8'b1101110;
DRAM[4005] = 8'b1101101;
DRAM[4006] = 8'b1101100;
DRAM[4007] = 8'b1101100;
DRAM[4008] = 8'b1101011;
DRAM[4009] = 8'b1101011;
DRAM[4010] = 8'b1101011;
DRAM[4011] = 8'b1101010;
DRAM[4012] = 8'b1101010;
DRAM[4013] = 8'b1101001;
DRAM[4014] = 8'b1101001;
DRAM[4015] = 8'b1101001;
DRAM[4016] = 8'b1101010;
DRAM[4017] = 8'b1101010;
DRAM[4018] = 8'b1101001;
DRAM[4019] = 8'b1101001;
DRAM[4020] = 8'b1101000;
DRAM[4021] = 8'b1100111;
DRAM[4022] = 8'b1100110;
DRAM[4023] = 8'b1100110;
DRAM[4024] = 8'b1100101;
DRAM[4025] = 8'b1100101;
DRAM[4026] = 8'b1100100;
DRAM[4027] = 8'b1100100;
DRAM[4028] = 8'b1100011;
DRAM[4029] = 8'b1100010;
DRAM[4030] = 8'b1100001;
DRAM[4031] = 8'b1100001;
DRAM[4032] = 8'b1100000;
DRAM[4033] = 8'b1100000;
DRAM[4034] = 8'b1011111;
DRAM[4035] = 8'b1011111;
DRAM[4036] = 8'b1011110;
DRAM[4037] = 8'b1011101;
DRAM[4038] = 8'b1011100;
DRAM[4039] = 8'b1011100;
DRAM[4040] = 8'b1011101;
DRAM[4041] = 8'b1011100;
DRAM[4042] = 8'b1011011;
DRAM[4043] = 8'b1011010;
DRAM[4044] = 8'b1011000;
DRAM[4045] = 8'b1010111;
DRAM[4046] = 8'b1010110;
DRAM[4047] = 8'b1010101;
DRAM[4048] = 8'b1010111;
DRAM[4049] = 8'b1010110;
DRAM[4050] = 8'b1010101;
DRAM[4051] = 8'b1010100;
DRAM[4052] = 8'b1010011;
DRAM[4053] = 8'b1010011;
DRAM[4054] = 8'b1010011;
DRAM[4055] = 8'b1010011;
DRAM[4056] = 8'b1001111;
DRAM[4057] = 8'b1001111;
DRAM[4058] = 8'b1001111;
DRAM[4059] = 8'b1001111;
DRAM[4060] = 8'b1001111;
DRAM[4061] = 8'b1001111;
DRAM[4062] = 8'b1001111;
DRAM[4063] = 8'b1001111;
DRAM[4064] = 8'b1001111;
DRAM[4065] = 8'b1001110;
DRAM[4066] = 8'b1001101;
DRAM[4067] = 8'b1001100;
DRAM[4068] = 8'b1001100;
DRAM[4069] = 8'b1001100;
DRAM[4070] = 8'b1001100;
DRAM[4071] = 8'b1001101;
DRAM[4072] = 8'b1001011;
DRAM[4073] = 8'b1001011;
DRAM[4074] = 8'b1001011;
DRAM[4075] = 8'b1001011;
DRAM[4076] = 8'b1001011;
DRAM[4077] = 8'b1001011;
DRAM[4078] = 8'b1001011;
DRAM[4079] = 8'b1001011;
DRAM[4080] = 8'b1001001;
DRAM[4081] = 8'b1001001;
DRAM[4082] = 8'b1001001;
DRAM[4083] = 8'b1001000;
DRAM[4084] = 8'b1001000;
DRAM[4085] = 8'b1001000;
DRAM[4086] = 8'b1000111;
DRAM[4087] = 8'b1000111;
DRAM[4088] = 8'b1000100;
DRAM[4089] = 8'b1000100;
DRAM[4090] = 8'b1000100;
DRAM[4091] = 8'b1000011;
DRAM[4092] = 8'b1000011;
DRAM[4093] = 8'b1000010;
DRAM[4094] = 8'b1000010;
DRAM[4095] = 8'b1000010;
DRAM[4096] = 8'b1100010;
DRAM[4097] = 8'b1100010;
DRAM[4098] = 8'b1100011;
DRAM[4099] = 8'b1100011;
DRAM[4100] = 8'b1100011;
DRAM[4101] = 8'b1100010;
DRAM[4102] = 8'b1100001;
DRAM[4103] = 8'b1100001;
DRAM[4104] = 8'b1100100;
DRAM[4105] = 8'b1100100;
DRAM[4106] = 8'b1100101;
DRAM[4107] = 8'b1100101;
DRAM[4108] = 8'b1100101;
DRAM[4109] = 8'b1100110;
DRAM[4110] = 8'b1100110;
DRAM[4111] = 8'b1100110;
DRAM[4112] = 8'b1100100;
DRAM[4113] = 8'b1100101;
DRAM[4114] = 8'b1100111;
DRAM[4115] = 8'b1101000;
DRAM[4116] = 8'b1101001;
DRAM[4117] = 8'b1101010;
DRAM[4118] = 8'b1101010;
DRAM[4119] = 8'b1101010;
DRAM[4120] = 8'b1101010;
DRAM[4121] = 8'b1101011;
DRAM[4122] = 8'b1101100;
DRAM[4123] = 8'b1101101;
DRAM[4124] = 8'b1101101;
DRAM[4125] = 8'b1101101;
DRAM[4126] = 8'b1101100;
DRAM[4127] = 8'b1101100;
DRAM[4128] = 8'b1101101;
DRAM[4129] = 8'b1101110;
DRAM[4130] = 8'b1101110;
DRAM[4131] = 8'b1101111;
DRAM[4132] = 8'b1101111;
DRAM[4133] = 8'b1101110;
DRAM[4134] = 8'b1101110;
DRAM[4135] = 8'b1101101;
DRAM[4136] = 8'b1101101;
DRAM[4137] = 8'b1101110;
DRAM[4138] = 8'b1101111;
DRAM[4139] = 8'b1101111;
DRAM[4140] = 8'b1110000;
DRAM[4141] = 8'b1110001;
DRAM[4142] = 8'b1110010;
DRAM[4143] = 8'b1110010;
DRAM[4144] = 8'b1110010;
DRAM[4145] = 8'b1110011;
DRAM[4146] = 8'b1110100;
DRAM[4147] = 8'b1110101;
DRAM[4148] = 8'b1110101;
DRAM[4149] = 8'b1110101;
DRAM[4150] = 8'b1110101;
DRAM[4151] = 8'b1110100;
DRAM[4152] = 8'b1110011;
DRAM[4153] = 8'b1110011;
DRAM[4154] = 8'b1110011;
DRAM[4155] = 8'b1110011;
DRAM[4156] = 8'b1110011;
DRAM[4157] = 8'b1110011;
DRAM[4158] = 8'b1110010;
DRAM[4159] = 8'b1110010;
DRAM[4160] = 8'b1110010;
DRAM[4161] = 8'b1110010;
DRAM[4162] = 8'b1110010;
DRAM[4163] = 8'b1110010;
DRAM[4164] = 8'b1110010;
DRAM[4165] = 8'b1110010;
DRAM[4166] = 8'b1110010;
DRAM[4167] = 8'b1110010;
DRAM[4168] = 8'b1110011;
DRAM[4169] = 8'b1110011;
DRAM[4170] = 8'b1110011;
DRAM[4171] = 8'b1110100;
DRAM[4172] = 8'b1110100;
DRAM[4173] = 8'b1110101;
DRAM[4174] = 8'b1110101;
DRAM[4175] = 8'b1110101;
DRAM[4176] = 8'b1110101;
DRAM[4177] = 8'b1110100;
DRAM[4178] = 8'b1110100;
DRAM[4179] = 8'b1110011;
DRAM[4180] = 8'b1110011;
DRAM[4181] = 8'b1110100;
DRAM[4182] = 8'b1110100;
DRAM[4183] = 8'b1110101;
DRAM[4184] = 8'b1110001;
DRAM[4185] = 8'b1110010;
DRAM[4186] = 8'b1110011;
DRAM[4187] = 8'b1110100;
DRAM[4188] = 8'b1110100;
DRAM[4189] = 8'b1110011;
DRAM[4190] = 8'b1110010;
DRAM[4191] = 8'b1110001;
DRAM[4192] = 8'b1110011;
DRAM[4193] = 8'b1110011;
DRAM[4194] = 8'b1110011;
DRAM[4195] = 8'b1110011;
DRAM[4196] = 8'b1110011;
DRAM[4197] = 8'b1110011;
DRAM[4198] = 8'b1110011;
DRAM[4199] = 8'b1110011;
DRAM[4200] = 8'b1110011;
DRAM[4201] = 8'b1110011;
DRAM[4202] = 8'b1110011;
DRAM[4203] = 8'b1110011;
DRAM[4204] = 8'b1110011;
DRAM[4205] = 8'b1110011;
DRAM[4206] = 8'b1110011;
DRAM[4207] = 8'b1110011;
DRAM[4208] = 8'b1110100;
DRAM[4209] = 8'b1110011;
DRAM[4210] = 8'b1110011;
DRAM[4211] = 8'b1110010;
DRAM[4212] = 8'b1110010;
DRAM[4213] = 8'b1110001;
DRAM[4214] = 8'b1110000;
DRAM[4215] = 8'b1110000;
DRAM[4216] = 8'b1110100;
DRAM[4217] = 8'b1110001;
DRAM[4218] = 8'b1101111;
DRAM[4219] = 8'b1110000;
DRAM[4220] = 8'b1110100;
DRAM[4221] = 8'b1110110;
DRAM[4222] = 8'b1110011;
DRAM[4223] = 8'b1110000;
DRAM[4224] = 8'b1110110;
DRAM[4225] = 8'b1110110;
DRAM[4226] = 8'b1110100;
DRAM[4227] = 8'b1110010;
DRAM[4228] = 8'b1101111;
DRAM[4229] = 8'b1101111;
DRAM[4230] = 8'b1110000;
DRAM[4231] = 8'b1110001;
DRAM[4232] = 8'b1110010;
DRAM[4233] = 8'b1110010;
DRAM[4234] = 8'b1110100;
DRAM[4235] = 8'b1110101;
DRAM[4236] = 8'b1110101;
DRAM[4237] = 8'b1110101;
DRAM[4238] = 8'b1110101;
DRAM[4239] = 8'b1110101;
DRAM[4240] = 8'b1110011;
DRAM[4241] = 8'b1110110;
DRAM[4242] = 8'b1110001;
DRAM[4243] = 8'b1110101;
DRAM[4244] = 8'b1110100;
DRAM[4245] = 8'b1110000;
DRAM[4246] = 8'b1110011;
DRAM[4247] = 8'b1101101;
DRAM[4248] = 8'b1110101;
DRAM[4249] = 8'b1110010;
DRAM[4250] = 8'b1110000;
DRAM[4251] = 8'b1110001;
DRAM[4252] = 8'b1110011;
DRAM[4253] = 8'b1110100;
DRAM[4254] = 8'b1110010;
DRAM[4255] = 8'b1110000;
DRAM[4256] = 8'b1110011;
DRAM[4257] = 8'b1101111;
DRAM[4258] = 8'b1101100;
DRAM[4259] = 8'b1101110;
DRAM[4260] = 8'b1110010;
DRAM[4261] = 8'b1110100;
DRAM[4262] = 8'b1110001;
DRAM[4263] = 8'b1101101;
DRAM[4264] = 8'b1101111;
DRAM[4265] = 8'b1101111;
DRAM[4266] = 8'b1101110;
DRAM[4267] = 8'b1101101;
DRAM[4268] = 8'b1101101;
DRAM[4269] = 8'b1101100;
DRAM[4270] = 8'b1101011;
DRAM[4271] = 8'b1101011;
DRAM[4272] = 8'b1101010;
DRAM[4273] = 8'b1101010;
DRAM[4274] = 8'b1101010;
DRAM[4275] = 8'b1101001;
DRAM[4276] = 8'b1101001;
DRAM[4277] = 8'b1101000;
DRAM[4278] = 8'b1101000;
DRAM[4279] = 8'b1101000;
DRAM[4280] = 8'b1100111;
DRAM[4281] = 8'b1100111;
DRAM[4282] = 8'b1100110;
DRAM[4283] = 8'b1100101;
DRAM[4284] = 8'b1100011;
DRAM[4285] = 8'b1100010;
DRAM[4286] = 8'b1100001;
DRAM[4287] = 8'b1100001;
DRAM[4288] = 8'b1100000;
DRAM[4289] = 8'b1100000;
DRAM[4290] = 8'b1100000;
DRAM[4291] = 8'b1100000;
DRAM[4292] = 8'b1011111;
DRAM[4293] = 8'b1011110;
DRAM[4294] = 8'b1011101;
DRAM[4295] = 8'b1011100;
DRAM[4296] = 8'b1011011;
DRAM[4297] = 8'b1011011;
DRAM[4298] = 8'b1011010;
DRAM[4299] = 8'b1011001;
DRAM[4300] = 8'b1011000;
DRAM[4301] = 8'b1011000;
DRAM[4302] = 8'b1010111;
DRAM[4303] = 8'b1010111;
DRAM[4304] = 8'b1010111;
DRAM[4305] = 8'b1010110;
DRAM[4306] = 8'b1010101;
DRAM[4307] = 8'b1010100;
DRAM[4308] = 8'b1010100;
DRAM[4309] = 8'b1010100;
DRAM[4310] = 8'b1010100;
DRAM[4311] = 8'b1010101;
DRAM[4312] = 8'b1010001;
DRAM[4313] = 8'b1010001;
DRAM[4314] = 8'b1010001;
DRAM[4315] = 8'b1010000;
DRAM[4316] = 8'b1010000;
DRAM[4317] = 8'b1001111;
DRAM[4318] = 8'b1001111;
DRAM[4319] = 8'b1001111;
DRAM[4320] = 8'b1001101;
DRAM[4321] = 8'b1001101;
DRAM[4322] = 8'b1001100;
DRAM[4323] = 8'b1001100;
DRAM[4324] = 8'b1001100;
DRAM[4325] = 8'b1001011;
DRAM[4326] = 8'b1001011;
DRAM[4327] = 8'b1001011;
DRAM[4328] = 8'b1001100;
DRAM[4329] = 8'b1001100;
DRAM[4330] = 8'b1001100;
DRAM[4331] = 8'b1001011;
DRAM[4332] = 8'b1001011;
DRAM[4333] = 8'b1001010;
DRAM[4334] = 8'b1001010;
DRAM[4335] = 8'b1001010;
DRAM[4336] = 8'b1001001;
DRAM[4337] = 8'b1001001;
DRAM[4338] = 8'b1001001;
DRAM[4339] = 8'b1001000;
DRAM[4340] = 8'b1001000;
DRAM[4341] = 8'b1000111;
DRAM[4342] = 8'b1000111;
DRAM[4343] = 8'b1000111;
DRAM[4344] = 8'b1000110;
DRAM[4345] = 8'b1000111;
DRAM[4346] = 8'b1000111;
DRAM[4347] = 8'b1000111;
DRAM[4348] = 8'b1000111;
DRAM[4349] = 8'b1000110;
DRAM[4350] = 8'b1000101;
DRAM[4351] = 8'b1000100;
DRAM[4352] = 8'b1100001;
DRAM[4353] = 8'b1100010;
DRAM[4354] = 8'b1100011;
DRAM[4355] = 8'b1100011;
DRAM[4356] = 8'b1100011;
DRAM[4357] = 8'b1100010;
DRAM[4358] = 8'b1100010;
DRAM[4359] = 8'b1100001;
DRAM[4360] = 8'b1100011;
DRAM[4361] = 8'b1100011;
DRAM[4362] = 8'b1100100;
DRAM[4363] = 8'b1100100;
DRAM[4364] = 8'b1100101;
DRAM[4365] = 8'b1100110;
DRAM[4366] = 8'b1100110;
DRAM[4367] = 8'b1100110;
DRAM[4368] = 8'b1100100;
DRAM[4369] = 8'b1100101;
DRAM[4370] = 8'b1100111;
DRAM[4371] = 8'b1101000;
DRAM[4372] = 8'b1101010;
DRAM[4373] = 8'b1101010;
DRAM[4374] = 8'b1101010;
DRAM[4375] = 8'b1101010;
DRAM[4376] = 8'b1101010;
DRAM[4377] = 8'b1101011;
DRAM[4378] = 8'b1101100;
DRAM[4379] = 8'b1101101;
DRAM[4380] = 8'b1101101;
DRAM[4381] = 8'b1101101;
DRAM[4382] = 8'b1101101;
DRAM[4383] = 8'b1101100;
DRAM[4384] = 8'b1101101;
DRAM[4385] = 8'b1101110;
DRAM[4386] = 8'b1101111;
DRAM[4387] = 8'b1101111;
DRAM[4388] = 8'b1101111;
DRAM[4389] = 8'b1101111;
DRAM[4390] = 8'b1101110;
DRAM[4391] = 8'b1101101;
DRAM[4392] = 8'b1101110;
DRAM[4393] = 8'b1101110;
DRAM[4394] = 8'b1101111;
DRAM[4395] = 8'b1110000;
DRAM[4396] = 8'b1110001;
DRAM[4397] = 8'b1110001;
DRAM[4398] = 8'b1110010;
DRAM[4399] = 8'b1110010;
DRAM[4400] = 8'b1110010;
DRAM[4401] = 8'b1110011;
DRAM[4402] = 8'b1110100;
DRAM[4403] = 8'b1110101;
DRAM[4404] = 8'b1110101;
DRAM[4405] = 8'b1110101;
DRAM[4406] = 8'b1110101;
DRAM[4407] = 8'b1110100;
DRAM[4408] = 8'b1110100;
DRAM[4409] = 8'b1110100;
DRAM[4410] = 8'b1110100;
DRAM[4411] = 8'b1110100;
DRAM[4412] = 8'b1110100;
DRAM[4413] = 8'b1110100;
DRAM[4414] = 8'b1110100;
DRAM[4415] = 8'b1110011;
DRAM[4416] = 8'b1110010;
DRAM[4417] = 8'b1110010;
DRAM[4418] = 8'b1110010;
DRAM[4419] = 8'b1110010;
DRAM[4420] = 8'b1110010;
DRAM[4421] = 8'b1110010;
DRAM[4422] = 8'b1110010;
DRAM[4423] = 8'b1110010;
DRAM[4424] = 8'b1110100;
DRAM[4425] = 8'b1110100;
DRAM[4426] = 8'b1110100;
DRAM[4427] = 8'b1110101;
DRAM[4428] = 8'b1110101;
DRAM[4429] = 8'b1110110;
DRAM[4430] = 8'b1110110;
DRAM[4431] = 8'b1110110;
DRAM[4432] = 8'b1110101;
DRAM[4433] = 8'b1110100;
DRAM[4434] = 8'b1110100;
DRAM[4435] = 8'b1110011;
DRAM[4436] = 8'b1110011;
DRAM[4437] = 8'b1110100;
DRAM[4438] = 8'b1110100;
DRAM[4439] = 8'b1110101;
DRAM[4440] = 8'b1110010;
DRAM[4441] = 8'b1110011;
DRAM[4442] = 8'b1110100;
DRAM[4443] = 8'b1110101;
DRAM[4444] = 8'b1110101;
DRAM[4445] = 8'b1110100;
DRAM[4446] = 8'b1110011;
DRAM[4447] = 8'b1110010;
DRAM[4448] = 8'b1110011;
DRAM[4449] = 8'b1110011;
DRAM[4450] = 8'b1110011;
DRAM[4451] = 8'b1110011;
DRAM[4452] = 8'b1110011;
DRAM[4453] = 8'b1110011;
DRAM[4454] = 8'b1110011;
DRAM[4455] = 8'b1110011;
DRAM[4456] = 8'b1110011;
DRAM[4457] = 8'b1110011;
DRAM[4458] = 8'b1110011;
DRAM[4459] = 8'b1110011;
DRAM[4460] = 8'b1110011;
DRAM[4461] = 8'b1110011;
DRAM[4462] = 8'b1110011;
DRAM[4463] = 8'b1110011;
DRAM[4464] = 8'b1110011;
DRAM[4465] = 8'b1110011;
DRAM[4466] = 8'b1110011;
DRAM[4467] = 8'b1110011;
DRAM[4468] = 8'b1110011;
DRAM[4469] = 8'b1110100;
DRAM[4470] = 8'b1110100;
DRAM[4471] = 8'b1110100;
DRAM[4472] = 8'b1110010;
DRAM[4473] = 8'b1110011;
DRAM[4474] = 8'b1110100;
DRAM[4475] = 8'b1110011;
DRAM[4476] = 8'b1110010;
DRAM[4477] = 8'b1110010;
DRAM[4478] = 8'b1110011;
DRAM[4479] = 8'b1110011;
DRAM[4480] = 8'b1110001;
DRAM[4481] = 8'b1110010;
DRAM[4482] = 8'b1110100;
DRAM[4483] = 8'b1110101;
DRAM[4484] = 8'b1110100;
DRAM[4485] = 8'b1110011;
DRAM[4486] = 8'b1110011;
DRAM[4487] = 8'b1110011;
DRAM[4488] = 8'b1110001;
DRAM[4489] = 8'b1110001;
DRAM[4490] = 8'b1110010;
DRAM[4491] = 8'b1110011;
DRAM[4492] = 8'b1110011;
DRAM[4493] = 8'b1110011;
DRAM[4494] = 8'b1110100;
DRAM[4495] = 8'b1110100;
DRAM[4496] = 8'b1110000;
DRAM[4497] = 8'b1110000;
DRAM[4498] = 8'b1101101;
DRAM[4499] = 8'b1110000;
DRAM[4500] = 8'b1110011;
DRAM[4501] = 8'b1110011;
DRAM[4502] = 8'b1110110;
DRAM[4503] = 8'b1110010;
DRAM[4504] = 8'b1110101;
DRAM[4505] = 8'b1110011;
DRAM[4506] = 8'b1110010;
DRAM[4507] = 8'b1110011;
DRAM[4508] = 8'b1110101;
DRAM[4509] = 8'b1110101;
DRAM[4510] = 8'b1110011;
DRAM[4511] = 8'b1110001;
DRAM[4512] = 8'b1110010;
DRAM[4513] = 8'b1101111;
DRAM[4514] = 8'b1101101;
DRAM[4515] = 8'b1101110;
DRAM[4516] = 8'b1110001;
DRAM[4517] = 8'b1110010;
DRAM[4518] = 8'b1110000;
DRAM[4519] = 8'b1101110;
DRAM[4520] = 8'b1101111;
DRAM[4521] = 8'b1101111;
DRAM[4522] = 8'b1101110;
DRAM[4523] = 8'b1101110;
DRAM[4524] = 8'b1101101;
DRAM[4525] = 8'b1101100;
DRAM[4526] = 8'b1101011;
DRAM[4527] = 8'b1101011;
DRAM[4528] = 8'b1101010;
DRAM[4529] = 8'b1101010;
DRAM[4530] = 8'b1101010;
DRAM[4531] = 8'b1101001;
DRAM[4532] = 8'b1101001;
DRAM[4533] = 8'b1101001;
DRAM[4534] = 8'b1101000;
DRAM[4535] = 8'b1101000;
DRAM[4536] = 8'b1100111;
DRAM[4537] = 8'b1100111;
DRAM[4538] = 8'b1100110;
DRAM[4539] = 8'b1100101;
DRAM[4540] = 8'b1100100;
DRAM[4541] = 8'b1100010;
DRAM[4542] = 8'b1100001;
DRAM[4543] = 8'b1100001;
DRAM[4544] = 8'b1100000;
DRAM[4545] = 8'b1100001;
DRAM[4546] = 8'b1100001;
DRAM[4547] = 8'b1100000;
DRAM[4548] = 8'b1100000;
DRAM[4549] = 8'b1011110;
DRAM[4550] = 8'b1011101;
DRAM[4551] = 8'b1011100;
DRAM[4552] = 8'b1011011;
DRAM[4553] = 8'b1011011;
DRAM[4554] = 8'b1011010;
DRAM[4555] = 8'b1011010;
DRAM[4556] = 8'b1011001;
DRAM[4557] = 8'b1011000;
DRAM[4558] = 8'b1010111;
DRAM[4559] = 8'b1010111;
DRAM[4560] = 8'b1010111;
DRAM[4561] = 8'b1010110;
DRAM[4562] = 8'b1010101;
DRAM[4563] = 8'b1010101;
DRAM[4564] = 8'b1010100;
DRAM[4565] = 8'b1010100;
DRAM[4566] = 8'b1010101;
DRAM[4567] = 8'b1010101;
DRAM[4568] = 8'b1010010;
DRAM[4569] = 8'b1010010;
DRAM[4570] = 8'b1010010;
DRAM[4571] = 8'b1010010;
DRAM[4572] = 8'b1010001;
DRAM[4573] = 8'b1010001;
DRAM[4574] = 8'b1010000;
DRAM[4575] = 8'b1010000;
DRAM[4576] = 8'b1001101;
DRAM[4577] = 8'b1001101;
DRAM[4578] = 8'b1001101;
DRAM[4579] = 8'b1001100;
DRAM[4580] = 8'b1001100;
DRAM[4581] = 8'b1001100;
DRAM[4582] = 8'b1001011;
DRAM[4583] = 8'b1001011;
DRAM[4584] = 8'b1001100;
DRAM[4585] = 8'b1001100;
DRAM[4586] = 8'b1001100;
DRAM[4587] = 8'b1001011;
DRAM[4588] = 8'b1001011;
DRAM[4589] = 8'b1001011;
DRAM[4590] = 8'b1001010;
DRAM[4591] = 8'b1001010;
DRAM[4592] = 8'b1001001;
DRAM[4593] = 8'b1001001;
DRAM[4594] = 8'b1001001;
DRAM[4595] = 8'b1001000;
DRAM[4596] = 8'b1001000;
DRAM[4597] = 8'b1001000;
DRAM[4598] = 8'b1000111;
DRAM[4599] = 8'b1000111;
DRAM[4600] = 8'b1000110;
DRAM[4601] = 8'b1000111;
DRAM[4602] = 8'b1000111;
DRAM[4603] = 8'b1000111;
DRAM[4604] = 8'b1000111;
DRAM[4605] = 8'b1000110;
DRAM[4606] = 8'b1000101;
DRAM[4607] = 8'b1000100;
DRAM[4608] = 8'b1100001;
DRAM[4609] = 8'b1100010;
DRAM[4610] = 8'b1100011;
DRAM[4611] = 8'b1100011;
DRAM[4612] = 8'b1100011;
DRAM[4613] = 8'b1100011;
DRAM[4614] = 8'b1100010;
DRAM[4615] = 8'b1100010;
DRAM[4616] = 8'b1100001;
DRAM[4617] = 8'b1100010;
DRAM[4618] = 8'b1100011;
DRAM[4619] = 8'b1100011;
DRAM[4620] = 8'b1100100;
DRAM[4621] = 8'b1100101;
DRAM[4622] = 8'b1100110;
DRAM[4623] = 8'b1100110;
DRAM[4624] = 8'b1100100;
DRAM[4625] = 8'b1100101;
DRAM[4626] = 8'b1100111;
DRAM[4627] = 8'b1101001;
DRAM[4628] = 8'b1101010;
DRAM[4629] = 8'b1101011;
DRAM[4630] = 8'b1101011;
DRAM[4631] = 8'b1101011;
DRAM[4632] = 8'b1101011;
DRAM[4633] = 8'b1101100;
DRAM[4634] = 8'b1101101;
DRAM[4635] = 8'b1101101;
DRAM[4636] = 8'b1101110;
DRAM[4637] = 8'b1101110;
DRAM[4638] = 8'b1101101;
DRAM[4639] = 8'b1101101;
DRAM[4640] = 8'b1101110;
DRAM[4641] = 8'b1101110;
DRAM[4642] = 8'b1101111;
DRAM[4643] = 8'b1110000;
DRAM[4644] = 8'b1110000;
DRAM[4645] = 8'b1101111;
DRAM[4646] = 8'b1101110;
DRAM[4647] = 8'b1101110;
DRAM[4648] = 8'b1101111;
DRAM[4649] = 8'b1101111;
DRAM[4650] = 8'b1101111;
DRAM[4651] = 8'b1110000;
DRAM[4652] = 8'b1110001;
DRAM[4653] = 8'b1110001;
DRAM[4654] = 8'b1110010;
DRAM[4655] = 8'b1110010;
DRAM[4656] = 8'b1110010;
DRAM[4657] = 8'b1110011;
DRAM[4658] = 8'b1110100;
DRAM[4659] = 8'b1110101;
DRAM[4660] = 8'b1110101;
DRAM[4661] = 8'b1110101;
DRAM[4662] = 8'b1110101;
DRAM[4663] = 8'b1110100;
DRAM[4664] = 8'b1110101;
DRAM[4665] = 8'b1110101;
DRAM[4666] = 8'b1110101;
DRAM[4667] = 8'b1110101;
DRAM[4668] = 8'b1110101;
DRAM[4669] = 8'b1110101;
DRAM[4670] = 8'b1110101;
DRAM[4671] = 8'b1110101;
DRAM[4672] = 8'b1110011;
DRAM[4673] = 8'b1110011;
DRAM[4674] = 8'b1110011;
DRAM[4675] = 8'b1110011;
DRAM[4676] = 8'b1110011;
DRAM[4677] = 8'b1110011;
DRAM[4678] = 8'b1110011;
DRAM[4679] = 8'b1110011;
DRAM[4680] = 8'b1110101;
DRAM[4681] = 8'b1110101;
DRAM[4682] = 8'b1110101;
DRAM[4683] = 8'b1110101;
DRAM[4684] = 8'b1110110;
DRAM[4685] = 8'b1110110;
DRAM[4686] = 8'b1110110;
DRAM[4687] = 8'b1110110;
DRAM[4688] = 8'b1110101;
DRAM[4689] = 8'b1110101;
DRAM[4690] = 8'b1110100;
DRAM[4691] = 8'b1110100;
DRAM[4692] = 8'b1110100;
DRAM[4693] = 8'b1110100;
DRAM[4694] = 8'b1110101;
DRAM[4695] = 8'b1110101;
DRAM[4696] = 8'b1110100;
DRAM[4697] = 8'b1110101;
DRAM[4698] = 8'b1110101;
DRAM[4699] = 8'b1110110;
DRAM[4700] = 8'b1110110;
DRAM[4701] = 8'b1110101;
DRAM[4702] = 8'b1110101;
DRAM[4703] = 8'b1110100;
DRAM[4704] = 8'b1110100;
DRAM[4705] = 8'b1110100;
DRAM[4706] = 8'b1110100;
DRAM[4707] = 8'b1110100;
DRAM[4708] = 8'b1110100;
DRAM[4709] = 8'b1110100;
DRAM[4710] = 8'b1110100;
DRAM[4711] = 8'b1110100;
DRAM[4712] = 8'b1110100;
DRAM[4713] = 8'b1110100;
DRAM[4714] = 8'b1110100;
DRAM[4715] = 8'b1110100;
DRAM[4716] = 8'b1110100;
DRAM[4717] = 8'b1110100;
DRAM[4718] = 8'b1110100;
DRAM[4719] = 8'b1110100;
DRAM[4720] = 8'b1110010;
DRAM[4721] = 8'b1110011;
DRAM[4722] = 8'b1110011;
DRAM[4723] = 8'b1110100;
DRAM[4724] = 8'b1110101;
DRAM[4725] = 8'b1110110;
DRAM[4726] = 8'b1110110;
DRAM[4727] = 8'b1110111;
DRAM[4728] = 8'b1101101;
DRAM[4729] = 8'b1110001;
DRAM[4730] = 8'b1110101;
DRAM[4731] = 8'b1110100;
DRAM[4732] = 8'b1110000;
DRAM[4733] = 8'b1101111;
DRAM[4734] = 8'b1110010;
DRAM[4735] = 8'b1110110;
DRAM[4736] = 8'b1110000;
DRAM[4737] = 8'b1110010;
DRAM[4738] = 8'b1110101;
DRAM[4739] = 8'b1110111;
DRAM[4740] = 8'b1111000;
DRAM[4741] = 8'b1110110;
DRAM[4742] = 8'b1110100;
DRAM[4743] = 8'b1110010;
DRAM[4744] = 8'b1110001;
DRAM[4745] = 8'b1110001;
DRAM[4746] = 8'b1110001;
DRAM[4747] = 8'b1110001;
DRAM[4748] = 8'b1110001;
DRAM[4749] = 8'b1110010;
DRAM[4750] = 8'b1110011;
DRAM[4751] = 8'b1110011;
DRAM[4752] = 8'b1110101;
DRAM[4753] = 8'b1110001;
DRAM[4754] = 8'b1101111;
DRAM[4755] = 8'b1101110;
DRAM[4756] = 8'b1110000;
DRAM[4757] = 8'b1110010;
DRAM[4758] = 8'b1101111;
DRAM[4759] = 8'b1101101;
DRAM[4760] = 8'b1110001;
DRAM[4761] = 8'b1110000;
DRAM[4762] = 8'b1110000;
DRAM[4763] = 8'b1110001;
DRAM[4764] = 8'b1110010;
DRAM[4765] = 8'b1110010;
DRAM[4766] = 8'b1110001;
DRAM[4767] = 8'b1101111;
DRAM[4768] = 8'b1110000;
DRAM[4769] = 8'b1101111;
DRAM[4770] = 8'b1101111;
DRAM[4771] = 8'b1101111;
DRAM[4772] = 8'b1101111;
DRAM[4773] = 8'b1101111;
DRAM[4774] = 8'b1101111;
DRAM[4775] = 8'b1101111;
DRAM[4776] = 8'b1101111;
DRAM[4777] = 8'b1101111;
DRAM[4778] = 8'b1101111;
DRAM[4779] = 8'b1101110;
DRAM[4780] = 8'b1101101;
DRAM[4781] = 8'b1101100;
DRAM[4782] = 8'b1101100;
DRAM[4783] = 8'b1101011;
DRAM[4784] = 8'b1101010;
DRAM[4785] = 8'b1101010;
DRAM[4786] = 8'b1101010;
DRAM[4787] = 8'b1101010;
DRAM[4788] = 8'b1101001;
DRAM[4789] = 8'b1101001;
DRAM[4790] = 8'b1101001;
DRAM[4791] = 8'b1101000;
DRAM[4792] = 8'b1101000;
DRAM[4793] = 8'b1100111;
DRAM[4794] = 8'b1100110;
DRAM[4795] = 8'b1100101;
DRAM[4796] = 8'b1100100;
DRAM[4797] = 8'b1100011;
DRAM[4798] = 8'b1100010;
DRAM[4799] = 8'b1100001;
DRAM[4800] = 8'b1100001;
DRAM[4801] = 8'b1100001;
DRAM[4802] = 8'b1100001;
DRAM[4803] = 8'b1100001;
DRAM[4804] = 8'b1100000;
DRAM[4805] = 8'b1011111;
DRAM[4806] = 8'b1011101;
DRAM[4807] = 8'b1011101;
DRAM[4808] = 8'b1011100;
DRAM[4809] = 8'b1011100;
DRAM[4810] = 8'b1011011;
DRAM[4811] = 8'b1011010;
DRAM[4812] = 8'b1011001;
DRAM[4813] = 8'b1011001;
DRAM[4814] = 8'b1011000;
DRAM[4815] = 8'b1011000;
DRAM[4816] = 8'b1010111;
DRAM[4817] = 8'b1010111;
DRAM[4818] = 8'b1010110;
DRAM[4819] = 8'b1010101;
DRAM[4820] = 8'b1010100;
DRAM[4821] = 8'b1010100;
DRAM[4822] = 8'b1010101;
DRAM[4823] = 8'b1010101;
DRAM[4824] = 8'b1010100;
DRAM[4825] = 8'b1010100;
DRAM[4826] = 8'b1010011;
DRAM[4827] = 8'b1010011;
DRAM[4828] = 8'b1010010;
DRAM[4829] = 8'b1010010;
DRAM[4830] = 8'b1010010;
DRAM[4831] = 8'b1010010;
DRAM[4832] = 8'b1001110;
DRAM[4833] = 8'b1001110;
DRAM[4834] = 8'b1001101;
DRAM[4835] = 8'b1001101;
DRAM[4836] = 8'b1001101;
DRAM[4837] = 8'b1001100;
DRAM[4838] = 8'b1001100;
DRAM[4839] = 8'b1001100;
DRAM[4840] = 8'b1001100;
DRAM[4841] = 8'b1001100;
DRAM[4842] = 8'b1001100;
DRAM[4843] = 8'b1001100;
DRAM[4844] = 8'b1001011;
DRAM[4845] = 8'b1001011;
DRAM[4846] = 8'b1001011;
DRAM[4847] = 8'b1001010;
DRAM[4848] = 8'b1001001;
DRAM[4849] = 8'b1001001;
DRAM[4850] = 8'b1001001;
DRAM[4851] = 8'b1001001;
DRAM[4852] = 8'b1001000;
DRAM[4853] = 8'b1001000;
DRAM[4854] = 8'b1001000;
DRAM[4855] = 8'b1000111;
DRAM[4856] = 8'b1000111;
DRAM[4857] = 8'b1000111;
DRAM[4858] = 8'b1000111;
DRAM[4859] = 8'b1000111;
DRAM[4860] = 8'b1000111;
DRAM[4861] = 8'b1000110;
DRAM[4862] = 8'b1000101;
DRAM[4863] = 8'b1000101;
DRAM[4864] = 8'b1100001;
DRAM[4865] = 8'b1100010;
DRAM[4866] = 8'b1100011;
DRAM[4867] = 8'b1100011;
DRAM[4868] = 8'b1100100;
DRAM[4869] = 8'b1100100;
DRAM[4870] = 8'b1100011;
DRAM[4871] = 8'b1100011;
DRAM[4872] = 8'b1100001;
DRAM[4873] = 8'b1100001;
DRAM[4874] = 8'b1100010;
DRAM[4875] = 8'b1100011;
DRAM[4876] = 8'b1100100;
DRAM[4877] = 8'b1100101;
DRAM[4878] = 8'b1100110;
DRAM[4879] = 8'b1100111;
DRAM[4880] = 8'b1100101;
DRAM[4881] = 8'b1100110;
DRAM[4882] = 8'b1100111;
DRAM[4883] = 8'b1101001;
DRAM[4884] = 8'b1101010;
DRAM[4885] = 8'b1101011;
DRAM[4886] = 8'b1101011;
DRAM[4887] = 8'b1101011;
DRAM[4888] = 8'b1101100;
DRAM[4889] = 8'b1101100;
DRAM[4890] = 8'b1101101;
DRAM[4891] = 8'b1101110;
DRAM[4892] = 8'b1101111;
DRAM[4893] = 8'b1101111;
DRAM[4894] = 8'b1101110;
DRAM[4895] = 8'b1101110;
DRAM[4896] = 8'b1101111;
DRAM[4897] = 8'b1101111;
DRAM[4898] = 8'b1110000;
DRAM[4899] = 8'b1110000;
DRAM[4900] = 8'b1110000;
DRAM[4901] = 8'b1110000;
DRAM[4902] = 8'b1101111;
DRAM[4903] = 8'b1101111;
DRAM[4904] = 8'b1101111;
DRAM[4905] = 8'b1110000;
DRAM[4906] = 8'b1110000;
DRAM[4907] = 8'b1110001;
DRAM[4908] = 8'b1110001;
DRAM[4909] = 8'b1110010;
DRAM[4910] = 8'b1110010;
DRAM[4911] = 8'b1110010;
DRAM[4912] = 8'b1110010;
DRAM[4913] = 8'b1110011;
DRAM[4914] = 8'b1110100;
DRAM[4915] = 8'b1110101;
DRAM[4916] = 8'b1110101;
DRAM[4917] = 8'b1110101;
DRAM[4918] = 8'b1110101;
DRAM[4919] = 8'b1110100;
DRAM[4920] = 8'b1110101;
DRAM[4921] = 8'b1110101;
DRAM[4922] = 8'b1110110;
DRAM[4923] = 8'b1110110;
DRAM[4924] = 8'b1110110;
DRAM[4925] = 8'b1110110;
DRAM[4926] = 8'b1110111;
DRAM[4927] = 8'b1110111;
DRAM[4928] = 8'b1110100;
DRAM[4929] = 8'b1110100;
DRAM[4930] = 8'b1110100;
DRAM[4931] = 8'b1110100;
DRAM[4932] = 8'b1110100;
DRAM[4933] = 8'b1110100;
DRAM[4934] = 8'b1110100;
DRAM[4935] = 8'b1110100;
DRAM[4936] = 8'b1110101;
DRAM[4937] = 8'b1110101;
DRAM[4938] = 8'b1110101;
DRAM[4939] = 8'b1110101;
DRAM[4940] = 8'b1110101;
DRAM[4941] = 8'b1110101;
DRAM[4942] = 8'b1110101;
DRAM[4943] = 8'b1110101;
DRAM[4944] = 8'b1110110;
DRAM[4945] = 8'b1110101;
DRAM[4946] = 8'b1110100;
DRAM[4947] = 8'b1110100;
DRAM[4948] = 8'b1110100;
DRAM[4949] = 8'b1110100;
DRAM[4950] = 8'b1110101;
DRAM[4951] = 8'b1110110;
DRAM[4952] = 8'b1110110;
DRAM[4953] = 8'b1110110;
DRAM[4954] = 8'b1110110;
DRAM[4955] = 8'b1110110;
DRAM[4956] = 8'b1110110;
DRAM[4957] = 8'b1110110;
DRAM[4958] = 8'b1110110;
DRAM[4959] = 8'b1110110;
DRAM[4960] = 8'b1110101;
DRAM[4961] = 8'b1110101;
DRAM[4962] = 8'b1110101;
DRAM[4963] = 8'b1110101;
DRAM[4964] = 8'b1110101;
DRAM[4965] = 8'b1110101;
DRAM[4966] = 8'b1110101;
DRAM[4967] = 8'b1110101;
DRAM[4968] = 8'b1110101;
DRAM[4969] = 8'b1110101;
DRAM[4970] = 8'b1110101;
DRAM[4971] = 8'b1110101;
DRAM[4972] = 8'b1110101;
DRAM[4973] = 8'b1110101;
DRAM[4974] = 8'b1110101;
DRAM[4975] = 8'b1110101;
DRAM[4976] = 8'b1110011;
DRAM[4977] = 8'b1110011;
DRAM[4978] = 8'b1110100;
DRAM[4979] = 8'b1110100;
DRAM[4980] = 8'b1110101;
DRAM[4981] = 8'b1110101;
DRAM[4982] = 8'b1110101;
DRAM[4983] = 8'b1110110;
DRAM[4984] = 8'b1110000;
DRAM[4985] = 8'b1110011;
DRAM[4986] = 8'b1110101;
DRAM[4987] = 8'b1110101;
DRAM[4988] = 8'b1110100;
DRAM[4989] = 8'b1110100;
DRAM[4990] = 8'b1110110;
DRAM[4991] = 8'b1111001;
DRAM[4992] = 8'b1110101;
DRAM[4993] = 8'b1110101;
DRAM[4994] = 8'b1110101;
DRAM[4995] = 8'b1110110;
DRAM[4996] = 8'b1110110;
DRAM[4997] = 8'b1110101;
DRAM[4998] = 8'b1110001;
DRAM[4999] = 8'b1101111;
DRAM[5000] = 8'b1110011;
DRAM[5001] = 8'b1110011;
DRAM[5002] = 8'b1110010;
DRAM[5003] = 8'b1110001;
DRAM[5004] = 8'b1110001;
DRAM[5005] = 8'b1110010;
DRAM[5006] = 8'b1110011;
DRAM[5007] = 8'b1110100;
DRAM[5008] = 8'b1111010;
DRAM[5009] = 8'b1110100;
DRAM[5010] = 8'b1110111;
DRAM[5011] = 8'b1110011;
DRAM[5012] = 8'b1110100;
DRAM[5013] = 8'b1111000;
DRAM[5014] = 8'b1101111;
DRAM[5015] = 8'b1110000;
DRAM[5016] = 8'b1110000;
DRAM[5017] = 8'b1110000;
DRAM[5018] = 8'b1110000;
DRAM[5019] = 8'b1110001;
DRAM[5020] = 8'b1110011;
DRAM[5021] = 8'b1110011;
DRAM[5022] = 8'b1110011;
DRAM[5023] = 8'b1110010;
DRAM[5024] = 8'b1101111;
DRAM[5025] = 8'b1110000;
DRAM[5026] = 8'b1110001;
DRAM[5027] = 8'b1110000;
DRAM[5028] = 8'b1101111;
DRAM[5029] = 8'b1101110;
DRAM[5030] = 8'b1101111;
DRAM[5031] = 8'b1110000;
DRAM[5032] = 8'b1110000;
DRAM[5033] = 8'b1110000;
DRAM[5034] = 8'b1101111;
DRAM[5035] = 8'b1101110;
DRAM[5036] = 8'b1101101;
DRAM[5037] = 8'b1101101;
DRAM[5038] = 8'b1101100;
DRAM[5039] = 8'b1101100;
DRAM[5040] = 8'b1101011;
DRAM[5041] = 8'b1101011;
DRAM[5042] = 8'b1101010;
DRAM[5043] = 8'b1101010;
DRAM[5044] = 8'b1101010;
DRAM[5045] = 8'b1101001;
DRAM[5046] = 8'b1101001;
DRAM[5047] = 8'b1101001;
DRAM[5048] = 8'b1101000;
DRAM[5049] = 8'b1100111;
DRAM[5050] = 8'b1100111;
DRAM[5051] = 8'b1100101;
DRAM[5052] = 8'b1100100;
DRAM[5053] = 8'b1100011;
DRAM[5054] = 8'b1100010;
DRAM[5055] = 8'b1100010;
DRAM[5056] = 8'b1100001;
DRAM[5057] = 8'b1100001;
DRAM[5058] = 8'b1100001;
DRAM[5059] = 8'b1100001;
DRAM[5060] = 8'b1100000;
DRAM[5061] = 8'b1011111;
DRAM[5062] = 8'b1011110;
DRAM[5063] = 8'b1011101;
DRAM[5064] = 8'b1011101;
DRAM[5065] = 8'b1011100;
DRAM[5066] = 8'b1011100;
DRAM[5067] = 8'b1011011;
DRAM[5068] = 8'b1011010;
DRAM[5069] = 8'b1011001;
DRAM[5070] = 8'b1011001;
DRAM[5071] = 8'b1011001;
DRAM[5072] = 8'b1011000;
DRAM[5073] = 8'b1010111;
DRAM[5074] = 8'b1010110;
DRAM[5075] = 8'b1010101;
DRAM[5076] = 8'b1010101;
DRAM[5077] = 8'b1010101;
DRAM[5078] = 8'b1010101;
DRAM[5079] = 8'b1010110;
DRAM[5080] = 8'b1010100;
DRAM[5081] = 8'b1010011;
DRAM[5082] = 8'b1010011;
DRAM[5083] = 8'b1010011;
DRAM[5084] = 8'b1010010;
DRAM[5085] = 8'b1010010;
DRAM[5086] = 8'b1010010;
DRAM[5087] = 8'b1010001;
DRAM[5088] = 8'b1001111;
DRAM[5089] = 8'b1001110;
DRAM[5090] = 8'b1001110;
DRAM[5091] = 8'b1001110;
DRAM[5092] = 8'b1001101;
DRAM[5093] = 8'b1001101;
DRAM[5094] = 8'b1001101;
DRAM[5095] = 8'b1001101;
DRAM[5096] = 8'b1001101;
DRAM[5097] = 8'b1001101;
DRAM[5098] = 8'b1001100;
DRAM[5099] = 8'b1001100;
DRAM[5100] = 8'b1001100;
DRAM[5101] = 8'b1001011;
DRAM[5102] = 8'b1001011;
DRAM[5103] = 8'b1001011;
DRAM[5104] = 8'b1001010;
DRAM[5105] = 8'b1001010;
DRAM[5106] = 8'b1001001;
DRAM[5107] = 8'b1001001;
DRAM[5108] = 8'b1001001;
DRAM[5109] = 8'b1001000;
DRAM[5110] = 8'b1001000;
DRAM[5111] = 8'b1001000;
DRAM[5112] = 8'b1000111;
DRAM[5113] = 8'b1000111;
DRAM[5114] = 8'b1001000;
DRAM[5115] = 8'b1001000;
DRAM[5116] = 8'b1000111;
DRAM[5117] = 8'b1000111;
DRAM[5118] = 8'b1000110;
DRAM[5119] = 8'b1000101;
DRAM[5120] = 8'b1100001;
DRAM[5121] = 8'b1100010;
DRAM[5122] = 8'b1100011;
DRAM[5123] = 8'b1100100;
DRAM[5124] = 8'b1100100;
DRAM[5125] = 8'b1100100;
DRAM[5126] = 8'b1100100;
DRAM[5127] = 8'b1100100;
DRAM[5128] = 8'b1100010;
DRAM[5129] = 8'b1100010;
DRAM[5130] = 8'b1100011;
DRAM[5131] = 8'b1100100;
DRAM[5132] = 8'b1100101;
DRAM[5133] = 8'b1100101;
DRAM[5134] = 8'b1100110;
DRAM[5135] = 8'b1100110;
DRAM[5136] = 8'b1100101;
DRAM[5137] = 8'b1100110;
DRAM[5138] = 8'b1101000;
DRAM[5139] = 8'b1101001;
DRAM[5140] = 8'b1101011;
DRAM[5141] = 8'b1101011;
DRAM[5142] = 8'b1101100;
DRAM[5143] = 8'b1101100;
DRAM[5144] = 8'b1101101;
DRAM[5145] = 8'b1101101;
DRAM[5146] = 8'b1101110;
DRAM[5147] = 8'b1101111;
DRAM[5148] = 8'b1101111;
DRAM[5149] = 8'b1101111;
DRAM[5150] = 8'b1101111;
DRAM[5151] = 8'b1101111;
DRAM[5152] = 8'b1110000;
DRAM[5153] = 8'b1110000;
DRAM[5154] = 8'b1110001;
DRAM[5155] = 8'b1110001;
DRAM[5156] = 8'b1110001;
DRAM[5157] = 8'b1110001;
DRAM[5158] = 8'b1110000;
DRAM[5159] = 8'b1110000;
DRAM[5160] = 8'b1110000;
DRAM[5161] = 8'b1110001;
DRAM[5162] = 8'b1110001;
DRAM[5163] = 8'b1110001;
DRAM[5164] = 8'b1110001;
DRAM[5165] = 8'b1110010;
DRAM[5166] = 8'b1110010;
DRAM[5167] = 8'b1110010;
DRAM[5168] = 8'b1110010;
DRAM[5169] = 8'b1110011;
DRAM[5170] = 8'b1110100;
DRAM[5171] = 8'b1110101;
DRAM[5172] = 8'b1110101;
DRAM[5173] = 8'b1110101;
DRAM[5174] = 8'b1110101;
DRAM[5175] = 8'b1110100;
DRAM[5176] = 8'b1110101;
DRAM[5177] = 8'b1110101;
DRAM[5178] = 8'b1110110;
DRAM[5179] = 8'b1110110;
DRAM[5180] = 8'b1110111;
DRAM[5181] = 8'b1110111;
DRAM[5182] = 8'b1110111;
DRAM[5183] = 8'b1111000;
DRAM[5184] = 8'b1110110;
DRAM[5185] = 8'b1110110;
DRAM[5186] = 8'b1110110;
DRAM[5187] = 8'b1110110;
DRAM[5188] = 8'b1110110;
DRAM[5189] = 8'b1110110;
DRAM[5190] = 8'b1110110;
DRAM[5191] = 8'b1110110;
DRAM[5192] = 8'b1110101;
DRAM[5193] = 8'b1110101;
DRAM[5194] = 8'b1110101;
DRAM[5195] = 8'b1110101;
DRAM[5196] = 8'b1110101;
DRAM[5197] = 8'b1110100;
DRAM[5198] = 8'b1110100;
DRAM[5199] = 8'b1110100;
DRAM[5200] = 8'b1110110;
DRAM[5201] = 8'b1110110;
DRAM[5202] = 8'b1110101;
DRAM[5203] = 8'b1110100;
DRAM[5204] = 8'b1110100;
DRAM[5205] = 8'b1110101;
DRAM[5206] = 8'b1110110;
DRAM[5207] = 8'b1110110;
DRAM[5208] = 8'b1110111;
DRAM[5209] = 8'b1110110;
DRAM[5210] = 8'b1110110;
DRAM[5211] = 8'b1110110;
DRAM[5212] = 8'b1110110;
DRAM[5213] = 8'b1110110;
DRAM[5214] = 8'b1110110;
DRAM[5215] = 8'b1110111;
DRAM[5216] = 8'b1110101;
DRAM[5217] = 8'b1110101;
DRAM[5218] = 8'b1110101;
DRAM[5219] = 8'b1110101;
DRAM[5220] = 8'b1110101;
DRAM[5221] = 8'b1110101;
DRAM[5222] = 8'b1110101;
DRAM[5223] = 8'b1110101;
DRAM[5224] = 8'b1110101;
DRAM[5225] = 8'b1110101;
DRAM[5226] = 8'b1110101;
DRAM[5227] = 8'b1110101;
DRAM[5228] = 8'b1110101;
DRAM[5229] = 8'b1110101;
DRAM[5230] = 8'b1110101;
DRAM[5231] = 8'b1110101;
DRAM[5232] = 8'b1110101;
DRAM[5233] = 8'b1110101;
DRAM[5234] = 8'b1110100;
DRAM[5235] = 8'b1110100;
DRAM[5236] = 8'b1110011;
DRAM[5237] = 8'b1110011;
DRAM[5238] = 8'b1110011;
DRAM[5239] = 8'b1110010;
DRAM[5240] = 8'b1111010;
DRAM[5241] = 8'b1111000;
DRAM[5242] = 8'b1110110;
DRAM[5243] = 8'b1110110;
DRAM[5244] = 8'b1111000;
DRAM[5245] = 8'b1111001;
DRAM[5246] = 8'b1110111;
DRAM[5247] = 8'b1110101;
DRAM[5248] = 8'b1111000;
DRAM[5249] = 8'b1110101;
DRAM[5250] = 8'b1110011;
DRAM[5251] = 8'b1110010;
DRAM[5252] = 8'b1110100;
DRAM[5253] = 8'b1110100;
DRAM[5254] = 8'b1110011;
DRAM[5255] = 8'b1110001;
DRAM[5256] = 8'b1110110;
DRAM[5257] = 8'b1110110;
DRAM[5258] = 8'b1110101;
DRAM[5259] = 8'b1110101;
DRAM[5260] = 8'b1110101;
DRAM[5261] = 8'b1110101;
DRAM[5262] = 8'b1110101;
DRAM[5263] = 8'b1110101;
DRAM[5264] = 8'b1110110;
DRAM[5265] = 8'b1101111;
DRAM[5266] = 8'b1111011;
DRAM[5267] = 8'b1110110;
DRAM[5268] = 8'b1110111;
DRAM[5269] = 8'b1111111;
DRAM[5270] = 8'b1110011;
DRAM[5271] = 8'b1111010;
DRAM[5272] = 8'b1110100;
DRAM[5273] = 8'b1110101;
DRAM[5274] = 8'b1110101;
DRAM[5275] = 8'b1110101;
DRAM[5276] = 8'b1110110;
DRAM[5277] = 8'b1110110;
DRAM[5278] = 8'b1111000;
DRAM[5279] = 8'b1111001;
DRAM[5280] = 8'b1110000;
DRAM[5281] = 8'b1110010;
DRAM[5282] = 8'b1110010;
DRAM[5283] = 8'b1110001;
DRAM[5284] = 8'b1101111;
DRAM[5285] = 8'b1101110;
DRAM[5286] = 8'b1101111;
DRAM[5287] = 8'b1110000;
DRAM[5288] = 8'b1110000;
DRAM[5289] = 8'b1110000;
DRAM[5290] = 8'b1101111;
DRAM[5291] = 8'b1101111;
DRAM[5292] = 8'b1101110;
DRAM[5293] = 8'b1101101;
DRAM[5294] = 8'b1101100;
DRAM[5295] = 8'b1101100;
DRAM[5296] = 8'b1101011;
DRAM[5297] = 8'b1101011;
DRAM[5298] = 8'b1101011;
DRAM[5299] = 8'b1101010;
DRAM[5300] = 8'b1101010;
DRAM[5301] = 8'b1101010;
DRAM[5302] = 8'b1101001;
DRAM[5303] = 8'b1101001;
DRAM[5304] = 8'b1101000;
DRAM[5305] = 8'b1101000;
DRAM[5306] = 8'b1100111;
DRAM[5307] = 8'b1100110;
DRAM[5308] = 8'b1100101;
DRAM[5309] = 8'b1100011;
DRAM[5310] = 8'b1100011;
DRAM[5311] = 8'b1100010;
DRAM[5312] = 8'b1100001;
DRAM[5313] = 8'b1100010;
DRAM[5314] = 8'b1100010;
DRAM[5315] = 8'b1100001;
DRAM[5316] = 8'b1100001;
DRAM[5317] = 8'b1011111;
DRAM[5318] = 8'b1011110;
DRAM[5319] = 8'b1011101;
DRAM[5320] = 8'b1011101;
DRAM[5321] = 8'b1011101;
DRAM[5322] = 8'b1011101;
DRAM[5323] = 8'b1011100;
DRAM[5324] = 8'b1011011;
DRAM[5325] = 8'b1011010;
DRAM[5326] = 8'b1011010;
DRAM[5327] = 8'b1011001;
DRAM[5328] = 8'b1011000;
DRAM[5329] = 8'b1010111;
DRAM[5330] = 8'b1010110;
DRAM[5331] = 8'b1010110;
DRAM[5332] = 8'b1010101;
DRAM[5333] = 8'b1010101;
DRAM[5334] = 8'b1010110;
DRAM[5335] = 8'b1010110;
DRAM[5336] = 8'b1010011;
DRAM[5337] = 8'b1010010;
DRAM[5338] = 8'b1010010;
DRAM[5339] = 8'b1010010;
DRAM[5340] = 8'b1010001;
DRAM[5341] = 8'b1010001;
DRAM[5342] = 8'b1010001;
DRAM[5343] = 8'b1010000;
DRAM[5344] = 8'b1001111;
DRAM[5345] = 8'b1001111;
DRAM[5346] = 8'b1001111;
DRAM[5347] = 8'b1001111;
DRAM[5348] = 8'b1001110;
DRAM[5349] = 8'b1001110;
DRAM[5350] = 8'b1001110;
DRAM[5351] = 8'b1001101;
DRAM[5352] = 8'b1001101;
DRAM[5353] = 8'b1001101;
DRAM[5354] = 8'b1001101;
DRAM[5355] = 8'b1001100;
DRAM[5356] = 8'b1001100;
DRAM[5357] = 8'b1001100;
DRAM[5358] = 8'b1001011;
DRAM[5359] = 8'b1001011;
DRAM[5360] = 8'b1001010;
DRAM[5361] = 8'b1001010;
DRAM[5362] = 8'b1001010;
DRAM[5363] = 8'b1001001;
DRAM[5364] = 8'b1001001;
DRAM[5365] = 8'b1001001;
DRAM[5366] = 8'b1001000;
DRAM[5367] = 8'b1001000;
DRAM[5368] = 8'b1000111;
DRAM[5369] = 8'b1001000;
DRAM[5370] = 8'b1001000;
DRAM[5371] = 8'b1001000;
DRAM[5372] = 8'b1001000;
DRAM[5373] = 8'b1000111;
DRAM[5374] = 8'b1000110;
DRAM[5375] = 8'b1000101;
DRAM[5376] = 8'b1100001;
DRAM[5377] = 8'b1100010;
DRAM[5378] = 8'b1100011;
DRAM[5379] = 8'b1100100;
DRAM[5380] = 8'b1100101;
DRAM[5381] = 8'b1100101;
DRAM[5382] = 8'b1100101;
DRAM[5383] = 8'b1100101;
DRAM[5384] = 8'b1100100;
DRAM[5385] = 8'b1100100;
DRAM[5386] = 8'b1100101;
DRAM[5387] = 8'b1100101;
DRAM[5388] = 8'b1100101;
DRAM[5389] = 8'b1100110;
DRAM[5390] = 8'b1100110;
DRAM[5391] = 8'b1100110;
DRAM[5392] = 8'b1100110;
DRAM[5393] = 8'b1100111;
DRAM[5394] = 8'b1101000;
DRAM[5395] = 8'b1101010;
DRAM[5396] = 8'b1101011;
DRAM[5397] = 8'b1101100;
DRAM[5398] = 8'b1101100;
DRAM[5399] = 8'b1101100;
DRAM[5400] = 8'b1101101;
DRAM[5401] = 8'b1101110;
DRAM[5402] = 8'b1101111;
DRAM[5403] = 8'b1110000;
DRAM[5404] = 8'b1110000;
DRAM[5405] = 8'b1110000;
DRAM[5406] = 8'b1110000;
DRAM[5407] = 8'b1101111;
DRAM[5408] = 8'b1110000;
DRAM[5409] = 8'b1110001;
DRAM[5410] = 8'b1110010;
DRAM[5411] = 8'b1110010;
DRAM[5412] = 8'b1110010;
DRAM[5413] = 8'b1110010;
DRAM[5414] = 8'b1110001;
DRAM[5415] = 8'b1110000;
DRAM[5416] = 8'b1110001;
DRAM[5417] = 8'b1110001;
DRAM[5418] = 8'b1110001;
DRAM[5419] = 8'b1110010;
DRAM[5420] = 8'b1110010;
DRAM[5421] = 8'b1110010;
DRAM[5422] = 8'b1110010;
DRAM[5423] = 8'b1110010;
DRAM[5424] = 8'b1110010;
DRAM[5425] = 8'b1110011;
DRAM[5426] = 8'b1110100;
DRAM[5427] = 8'b1110101;
DRAM[5428] = 8'b1110101;
DRAM[5429] = 8'b1110101;
DRAM[5430] = 8'b1110101;
DRAM[5431] = 8'b1110100;
DRAM[5432] = 8'b1110100;
DRAM[5433] = 8'b1110100;
DRAM[5434] = 8'b1110101;
DRAM[5435] = 8'b1110110;
DRAM[5436] = 8'b1110110;
DRAM[5437] = 8'b1110111;
DRAM[5438] = 8'b1111000;
DRAM[5439] = 8'b1111000;
DRAM[5440] = 8'b1110111;
DRAM[5441] = 8'b1110111;
DRAM[5442] = 8'b1110111;
DRAM[5443] = 8'b1110111;
DRAM[5444] = 8'b1110111;
DRAM[5445] = 8'b1110111;
DRAM[5446] = 8'b1110111;
DRAM[5447] = 8'b1110111;
DRAM[5448] = 8'b1110110;
DRAM[5449] = 8'b1110110;
DRAM[5450] = 8'b1110110;
DRAM[5451] = 8'b1110110;
DRAM[5452] = 8'b1110101;
DRAM[5453] = 8'b1110101;
DRAM[5454] = 8'b1110101;
DRAM[5455] = 8'b1110101;
DRAM[5456] = 8'b1110110;
DRAM[5457] = 8'b1110110;
DRAM[5458] = 8'b1110101;
DRAM[5459] = 8'b1110101;
DRAM[5460] = 8'b1110101;
DRAM[5461] = 8'b1110101;
DRAM[5462] = 8'b1110110;
DRAM[5463] = 8'b1110110;
DRAM[5464] = 8'b1110111;
DRAM[5465] = 8'b1110110;
DRAM[5466] = 8'b1110110;
DRAM[5467] = 8'b1110101;
DRAM[5468] = 8'b1110101;
DRAM[5469] = 8'b1110110;
DRAM[5470] = 8'b1110110;
DRAM[5471] = 8'b1110111;
DRAM[5472] = 8'b1110110;
DRAM[5473] = 8'b1110110;
DRAM[5474] = 8'b1110110;
DRAM[5475] = 8'b1110110;
DRAM[5476] = 8'b1110110;
DRAM[5477] = 8'b1110110;
DRAM[5478] = 8'b1110110;
DRAM[5479] = 8'b1110110;
DRAM[5480] = 8'b1110110;
DRAM[5481] = 8'b1110110;
DRAM[5482] = 8'b1110110;
DRAM[5483] = 8'b1110110;
DRAM[5484] = 8'b1110110;
DRAM[5485] = 8'b1110110;
DRAM[5486] = 8'b1110110;
DRAM[5487] = 8'b1110110;
DRAM[5488] = 8'b1110110;
DRAM[5489] = 8'b1110101;
DRAM[5490] = 8'b1110101;
DRAM[5491] = 8'b1110100;
DRAM[5492] = 8'b1110011;
DRAM[5493] = 8'b1110010;
DRAM[5494] = 8'b1110010;
DRAM[5495] = 8'b1110001;
DRAM[5496] = 8'b1111011;
DRAM[5497] = 8'b1110110;
DRAM[5498] = 8'b1110010;
DRAM[5499] = 8'b1110010;
DRAM[5500] = 8'b1110101;
DRAM[5501] = 8'b1110101;
DRAM[5502] = 8'b1110001;
DRAM[5503] = 8'b1101101;
DRAM[5504] = 8'b1110110;
DRAM[5505] = 8'b1110011;
DRAM[5506] = 8'b1110000;
DRAM[5507] = 8'b1110001;
DRAM[5508] = 8'b1110110;
DRAM[5509] = 8'b1111001;
DRAM[5510] = 8'b1111001;
DRAM[5511] = 8'b1110111;
DRAM[5512] = 8'b1110111;
DRAM[5513] = 8'b1111000;
DRAM[5514] = 8'b1111000;
DRAM[5515] = 8'b1111001;
DRAM[5516] = 8'b1111000;
DRAM[5517] = 8'b1110111;
DRAM[5518] = 8'b1110110;
DRAM[5519] = 8'b1110110;
DRAM[5520] = 8'b1110100;
DRAM[5521] = 8'b1101011;
DRAM[5522] = 8'b1111101;
DRAM[5523] = 8'b1110000;
DRAM[5524] = 8'b1101101;
DRAM[5525] = 8'b1111000;
DRAM[5526] = 8'b1101100;
DRAM[5527] = 8'b1111011;
DRAM[5528] = 8'b1111010;
DRAM[5529] = 8'b1111001;
DRAM[5530] = 8'b1111000;
DRAM[5531] = 8'b1110101;
DRAM[5532] = 8'b1110010;
DRAM[5533] = 8'b1110010;
DRAM[5534] = 8'b1110101;
DRAM[5535] = 8'b1111000;
DRAM[5536] = 8'b1110100;
DRAM[5537] = 8'b1110011;
DRAM[5538] = 8'b1110011;
DRAM[5539] = 8'b1110010;
DRAM[5540] = 8'b1110001;
DRAM[5541] = 8'b1110001;
DRAM[5542] = 8'b1110000;
DRAM[5543] = 8'b1110000;
DRAM[5544] = 8'b1110001;
DRAM[5545] = 8'b1110000;
DRAM[5546] = 8'b1110000;
DRAM[5547] = 8'b1101111;
DRAM[5548] = 8'b1101110;
DRAM[5549] = 8'b1101101;
DRAM[5550] = 8'b1101101;
DRAM[5551] = 8'b1101101;
DRAM[5552] = 8'b1101100;
DRAM[5553] = 8'b1101011;
DRAM[5554] = 8'b1101011;
DRAM[5555] = 8'b1101011;
DRAM[5556] = 8'b1101010;
DRAM[5557] = 8'b1101010;
DRAM[5558] = 8'b1101010;
DRAM[5559] = 8'b1101010;
DRAM[5560] = 8'b1101001;
DRAM[5561] = 8'b1101000;
DRAM[5562] = 8'b1100111;
DRAM[5563] = 8'b1100110;
DRAM[5564] = 8'b1100101;
DRAM[5565] = 8'b1100100;
DRAM[5566] = 8'b1100011;
DRAM[5567] = 8'b1100010;
DRAM[5568] = 8'b1100010;
DRAM[5569] = 8'b1100010;
DRAM[5570] = 8'b1100010;
DRAM[5571] = 8'b1100010;
DRAM[5572] = 8'b1100001;
DRAM[5573] = 8'b1100000;
DRAM[5574] = 8'b1011110;
DRAM[5575] = 8'b1011110;
DRAM[5576] = 8'b1011110;
DRAM[5577] = 8'b1011110;
DRAM[5578] = 8'b1011101;
DRAM[5579] = 8'b1011101;
DRAM[5580] = 8'b1011100;
DRAM[5581] = 8'b1011011;
DRAM[5582] = 8'b1011010;
DRAM[5583] = 8'b1011010;
DRAM[5584] = 8'b1011000;
DRAM[5585] = 8'b1011000;
DRAM[5586] = 8'b1010111;
DRAM[5587] = 8'b1010110;
DRAM[5588] = 8'b1010110;
DRAM[5589] = 8'b1010110;
DRAM[5590] = 8'b1010110;
DRAM[5591] = 8'b1010110;
DRAM[5592] = 8'b1010010;
DRAM[5593] = 8'b1010010;
DRAM[5594] = 8'b1010010;
DRAM[5595] = 8'b1010010;
DRAM[5596] = 8'b1010001;
DRAM[5597] = 8'b1010001;
DRAM[5598] = 8'b1010000;
DRAM[5599] = 8'b1010000;
DRAM[5600] = 8'b1010000;
DRAM[5601] = 8'b1010000;
DRAM[5602] = 8'b1010000;
DRAM[5603] = 8'b1001111;
DRAM[5604] = 8'b1001111;
DRAM[5605] = 8'b1001111;
DRAM[5606] = 8'b1001110;
DRAM[5607] = 8'b1001110;
DRAM[5608] = 8'b1001110;
DRAM[5609] = 8'b1001101;
DRAM[5610] = 8'b1001101;
DRAM[5611] = 8'b1001101;
DRAM[5612] = 8'b1001100;
DRAM[5613] = 8'b1001100;
DRAM[5614] = 8'b1001100;
DRAM[5615] = 8'b1001100;
DRAM[5616] = 8'b1001011;
DRAM[5617] = 8'b1001010;
DRAM[5618] = 8'b1001010;
DRAM[5619] = 8'b1001010;
DRAM[5620] = 8'b1001001;
DRAM[5621] = 8'b1001001;
DRAM[5622] = 8'b1001001;
DRAM[5623] = 8'b1001001;
DRAM[5624] = 8'b1001000;
DRAM[5625] = 8'b1001000;
DRAM[5626] = 8'b1001001;
DRAM[5627] = 8'b1001001;
DRAM[5628] = 8'b1001000;
DRAM[5629] = 8'b1000111;
DRAM[5630] = 8'b1000110;
DRAM[5631] = 8'b1000110;
DRAM[5632] = 8'b1100001;
DRAM[5633] = 8'b1100010;
DRAM[5634] = 8'b1100011;
DRAM[5635] = 8'b1100100;
DRAM[5636] = 8'b1100101;
DRAM[5637] = 8'b1100101;
DRAM[5638] = 8'b1100101;
DRAM[5639] = 8'b1100101;
DRAM[5640] = 8'b1100111;
DRAM[5641] = 8'b1100111;
DRAM[5642] = 8'b1100111;
DRAM[5643] = 8'b1100111;
DRAM[5644] = 8'b1100110;
DRAM[5645] = 8'b1100110;
DRAM[5646] = 8'b1100110;
DRAM[5647] = 8'b1100110;
DRAM[5648] = 8'b1100110;
DRAM[5649] = 8'b1100111;
DRAM[5650] = 8'b1101000;
DRAM[5651] = 8'b1101010;
DRAM[5652] = 8'b1101011;
DRAM[5653] = 8'b1101100;
DRAM[5654] = 8'b1101100;
DRAM[5655] = 8'b1101100;
DRAM[5656] = 8'b1101110;
DRAM[5657] = 8'b1101111;
DRAM[5658] = 8'b1101111;
DRAM[5659] = 8'b1110000;
DRAM[5660] = 8'b1110001;
DRAM[5661] = 8'b1110001;
DRAM[5662] = 8'b1110000;
DRAM[5663] = 8'b1110000;
DRAM[5664] = 8'b1110001;
DRAM[5665] = 8'b1110001;
DRAM[5666] = 8'b1110010;
DRAM[5667] = 8'b1110011;
DRAM[5668] = 8'b1110011;
DRAM[5669] = 8'b1110010;
DRAM[5670] = 8'b1110001;
DRAM[5671] = 8'b1110001;
DRAM[5672] = 8'b1110010;
DRAM[5673] = 8'b1110010;
DRAM[5674] = 8'b1110010;
DRAM[5675] = 8'b1110010;
DRAM[5676] = 8'b1110010;
DRAM[5677] = 8'b1110010;
DRAM[5678] = 8'b1110010;
DRAM[5679] = 8'b1110010;
DRAM[5680] = 8'b1110010;
DRAM[5681] = 8'b1110011;
DRAM[5682] = 8'b1110100;
DRAM[5683] = 8'b1110101;
DRAM[5684] = 8'b1110101;
DRAM[5685] = 8'b1110101;
DRAM[5686] = 8'b1110101;
DRAM[5687] = 8'b1110100;
DRAM[5688] = 8'b1110011;
DRAM[5689] = 8'b1110011;
DRAM[5690] = 8'b1110100;
DRAM[5691] = 8'b1110101;
DRAM[5692] = 8'b1110110;
DRAM[5693] = 8'b1110111;
DRAM[5694] = 8'b1110111;
DRAM[5695] = 8'b1111000;
DRAM[5696] = 8'b1111000;
DRAM[5697] = 8'b1111000;
DRAM[5698] = 8'b1111000;
DRAM[5699] = 8'b1111000;
DRAM[5700] = 8'b1111000;
DRAM[5701] = 8'b1111000;
DRAM[5702] = 8'b1111000;
DRAM[5703] = 8'b1111000;
DRAM[5704] = 8'b1111001;
DRAM[5705] = 8'b1111001;
DRAM[5706] = 8'b1111001;
DRAM[5707] = 8'b1111000;
DRAM[5708] = 8'b1111000;
DRAM[5709] = 8'b1110111;
DRAM[5710] = 8'b1110111;
DRAM[5711] = 8'b1110111;
DRAM[5712] = 8'b1110111;
DRAM[5713] = 8'b1110110;
DRAM[5714] = 8'b1110110;
DRAM[5715] = 8'b1110101;
DRAM[5716] = 8'b1110101;
DRAM[5717] = 8'b1110110;
DRAM[5718] = 8'b1110110;
DRAM[5719] = 8'b1110111;
DRAM[5720] = 8'b1110111;
DRAM[5721] = 8'b1110110;
DRAM[5722] = 8'b1110101;
DRAM[5723] = 8'b1110100;
DRAM[5724] = 8'b1110100;
DRAM[5725] = 8'b1110101;
DRAM[5726] = 8'b1110110;
DRAM[5727] = 8'b1110111;
DRAM[5728] = 8'b1110111;
DRAM[5729] = 8'b1110111;
DRAM[5730] = 8'b1110111;
DRAM[5731] = 8'b1110111;
DRAM[5732] = 8'b1110111;
DRAM[5733] = 8'b1110111;
DRAM[5734] = 8'b1110111;
DRAM[5735] = 8'b1110111;
DRAM[5736] = 8'b1110111;
DRAM[5737] = 8'b1110111;
DRAM[5738] = 8'b1110111;
DRAM[5739] = 8'b1110111;
DRAM[5740] = 8'b1110111;
DRAM[5741] = 8'b1110111;
DRAM[5742] = 8'b1110111;
DRAM[5743] = 8'b1110111;
DRAM[5744] = 8'b1110101;
DRAM[5745] = 8'b1110101;
DRAM[5746] = 8'b1110101;
DRAM[5747] = 8'b1110101;
DRAM[5748] = 8'b1110101;
DRAM[5749] = 8'b1110100;
DRAM[5750] = 8'b1110100;
DRAM[5751] = 8'b1110100;
DRAM[5752] = 8'b1110100;
DRAM[5753] = 8'b1110100;
DRAM[5754] = 8'b1110100;
DRAM[5755] = 8'b1110110;
DRAM[5756] = 8'b1111000;
DRAM[5757] = 8'b1111001;
DRAM[5758] = 8'b1111001;
DRAM[5759] = 8'b1111001;
DRAM[5760] = 8'b1110111;
DRAM[5761] = 8'b1110100;
DRAM[5762] = 8'b1110011;
DRAM[5763] = 8'b1110110;
DRAM[5764] = 8'b1111011;
DRAM[5765] = 8'b1111101;
DRAM[5766] = 8'b1111011;
DRAM[5767] = 8'b1111000;
DRAM[5768] = 8'b1110111;
DRAM[5769] = 8'b1111000;
DRAM[5770] = 8'b1111010;
DRAM[5771] = 8'b1111011;
DRAM[5772] = 8'b1111011;
DRAM[5773] = 8'b1111001;
DRAM[5774] = 8'b1110110;
DRAM[5775] = 8'b1110100;
DRAM[5776] = 8'b1111001;
DRAM[5777] = 8'b1101110;
DRAM[5778] = 8'b10000011;
DRAM[5779] = 8'b1110001;
DRAM[5780] = 8'b1101100;
DRAM[5781] = 8'b1111110;
DRAM[5782] = 8'b1110111;
DRAM[5783] = 8'b10010010;
DRAM[5784] = 8'b10000110;
DRAM[5785] = 8'b10000100;
DRAM[5786] = 8'b1111111;
DRAM[5787] = 8'b1110111;
DRAM[5788] = 8'b1110001;
DRAM[5789] = 8'b1110000;
DRAM[5790] = 8'b1110011;
DRAM[5791] = 8'b1110110;
DRAM[5792] = 8'b1111000;
DRAM[5793] = 8'b1110101;
DRAM[5794] = 8'b1110010;
DRAM[5795] = 8'b1110010;
DRAM[5796] = 8'b1110100;
DRAM[5797] = 8'b1110100;
DRAM[5798] = 8'b1110010;
DRAM[5799] = 8'b1101111;
DRAM[5800] = 8'b1110001;
DRAM[5801] = 8'b1110001;
DRAM[5802] = 8'b1110000;
DRAM[5803] = 8'b1101111;
DRAM[5804] = 8'b1101110;
DRAM[5805] = 8'b1101110;
DRAM[5806] = 8'b1101101;
DRAM[5807] = 8'b1101101;
DRAM[5808] = 8'b1101100;
DRAM[5809] = 8'b1101100;
DRAM[5810] = 8'b1101011;
DRAM[5811] = 8'b1101011;
DRAM[5812] = 8'b1101011;
DRAM[5813] = 8'b1101010;
DRAM[5814] = 8'b1101010;
DRAM[5815] = 8'b1101010;
DRAM[5816] = 8'b1101001;
DRAM[5817] = 8'b1101001;
DRAM[5818] = 8'b1101000;
DRAM[5819] = 8'b1100110;
DRAM[5820] = 8'b1100101;
DRAM[5821] = 8'b1100100;
DRAM[5822] = 8'b1100011;
DRAM[5823] = 8'b1100011;
DRAM[5824] = 8'b1100010;
DRAM[5825] = 8'b1100010;
DRAM[5826] = 8'b1100010;
DRAM[5827] = 8'b1100010;
DRAM[5828] = 8'b1100001;
DRAM[5829] = 8'b1100000;
DRAM[5830] = 8'b1011111;
DRAM[5831] = 8'b1011110;
DRAM[5832] = 8'b1011111;
DRAM[5833] = 8'b1011111;
DRAM[5834] = 8'b1011110;
DRAM[5835] = 8'b1011101;
DRAM[5836] = 8'b1011100;
DRAM[5837] = 8'b1011100;
DRAM[5838] = 8'b1011011;
DRAM[5839] = 8'b1011011;
DRAM[5840] = 8'b1011001;
DRAM[5841] = 8'b1011000;
DRAM[5842] = 8'b1010111;
DRAM[5843] = 8'b1010110;
DRAM[5844] = 8'b1010110;
DRAM[5845] = 8'b1010110;
DRAM[5846] = 8'b1010110;
DRAM[5847] = 8'b1010111;
DRAM[5848] = 8'b1010100;
DRAM[5849] = 8'b1010100;
DRAM[5850] = 8'b1010011;
DRAM[5851] = 8'b1010011;
DRAM[5852] = 8'b1010010;
DRAM[5853] = 8'b1010010;
DRAM[5854] = 8'b1010010;
DRAM[5855] = 8'b1010010;
DRAM[5856] = 8'b1010001;
DRAM[5857] = 8'b1010001;
DRAM[5858] = 8'b1010000;
DRAM[5859] = 8'b1010000;
DRAM[5860] = 8'b1010000;
DRAM[5861] = 8'b1001111;
DRAM[5862] = 8'b1001111;
DRAM[5863] = 8'b1001111;
DRAM[5864] = 8'b1001110;
DRAM[5865] = 8'b1001110;
DRAM[5866] = 8'b1001101;
DRAM[5867] = 8'b1001101;
DRAM[5868] = 8'b1001101;
DRAM[5869] = 8'b1001100;
DRAM[5870] = 8'b1001100;
DRAM[5871] = 8'b1001100;
DRAM[5872] = 8'b1001011;
DRAM[5873] = 8'b1001011;
DRAM[5874] = 8'b1001010;
DRAM[5875] = 8'b1001010;
DRAM[5876] = 8'b1001010;
DRAM[5877] = 8'b1001001;
DRAM[5878] = 8'b1001001;
DRAM[5879] = 8'b1001001;
DRAM[5880] = 8'b1001000;
DRAM[5881] = 8'b1001000;
DRAM[5882] = 8'b1001001;
DRAM[5883] = 8'b1001001;
DRAM[5884] = 8'b1001000;
DRAM[5885] = 8'b1001000;
DRAM[5886] = 8'b1000111;
DRAM[5887] = 8'b1000110;
DRAM[5888] = 8'b1100001;
DRAM[5889] = 8'b1100010;
DRAM[5890] = 8'b1100011;
DRAM[5891] = 8'b1100100;
DRAM[5892] = 8'b1100101;
DRAM[5893] = 8'b1100110;
DRAM[5894] = 8'b1100110;
DRAM[5895] = 8'b1100110;
DRAM[5896] = 8'b1101001;
DRAM[5897] = 8'b1101001;
DRAM[5898] = 8'b1101000;
DRAM[5899] = 8'b1101000;
DRAM[5900] = 8'b1100111;
DRAM[5901] = 8'b1100110;
DRAM[5902] = 8'b1100101;
DRAM[5903] = 8'b1100101;
DRAM[5904] = 8'b1100110;
DRAM[5905] = 8'b1100111;
DRAM[5906] = 8'b1101001;
DRAM[5907] = 8'b1101010;
DRAM[5908] = 8'b1101011;
DRAM[5909] = 8'b1101100;
DRAM[5910] = 8'b1101100;
DRAM[5911] = 8'b1101100;
DRAM[5912] = 8'b1101110;
DRAM[5913] = 8'b1101111;
DRAM[5914] = 8'b1110000;
DRAM[5915] = 8'b1110001;
DRAM[5916] = 8'b1110001;
DRAM[5917] = 8'b1110001;
DRAM[5918] = 8'b1110001;
DRAM[5919] = 8'b1110000;
DRAM[5920] = 8'b1110001;
DRAM[5921] = 8'b1110010;
DRAM[5922] = 8'b1110010;
DRAM[5923] = 8'b1110011;
DRAM[5924] = 8'b1110011;
DRAM[5925] = 8'b1110010;
DRAM[5926] = 8'b1110010;
DRAM[5927] = 8'b1110001;
DRAM[5928] = 8'b1110010;
DRAM[5929] = 8'b1110010;
DRAM[5930] = 8'b1110010;
DRAM[5931] = 8'b1110010;
DRAM[5932] = 8'b1110010;
DRAM[5933] = 8'b1110010;
DRAM[5934] = 8'b1110010;
DRAM[5935] = 8'b1110010;
DRAM[5936] = 8'b1110010;
DRAM[5937] = 8'b1110011;
DRAM[5938] = 8'b1110100;
DRAM[5939] = 8'b1110101;
DRAM[5940] = 8'b1110101;
DRAM[5941] = 8'b1110101;
DRAM[5942] = 8'b1110101;
DRAM[5943] = 8'b1110100;
DRAM[5944] = 8'b1110010;
DRAM[5945] = 8'b1110011;
DRAM[5946] = 8'b1110100;
DRAM[5947] = 8'b1110100;
DRAM[5948] = 8'b1110101;
DRAM[5949] = 8'b1110110;
DRAM[5950] = 8'b1110111;
DRAM[5951] = 8'b1110111;
DRAM[5952] = 8'b1111000;
DRAM[5953] = 8'b1111000;
DRAM[5954] = 8'b1111000;
DRAM[5955] = 8'b1111000;
DRAM[5956] = 8'b1111000;
DRAM[5957] = 8'b1111000;
DRAM[5958] = 8'b1111000;
DRAM[5959] = 8'b1111000;
DRAM[5960] = 8'b1111100;
DRAM[5961] = 8'b1111011;
DRAM[5962] = 8'b1111011;
DRAM[5963] = 8'b1111011;
DRAM[5964] = 8'b1111010;
DRAM[5965] = 8'b1111001;
DRAM[5966] = 8'b1111001;
DRAM[5967] = 8'b1111001;
DRAM[5968] = 8'b1110111;
DRAM[5969] = 8'b1110110;
DRAM[5970] = 8'b1110110;
DRAM[5971] = 8'b1110101;
DRAM[5972] = 8'b1110101;
DRAM[5973] = 8'b1110110;
DRAM[5974] = 8'b1110110;
DRAM[5975] = 8'b1110111;
DRAM[5976] = 8'b1110110;
DRAM[5977] = 8'b1110110;
DRAM[5978] = 8'b1110100;
DRAM[5979] = 8'b1110011;
DRAM[5980] = 8'b1110011;
DRAM[5981] = 8'b1110100;
DRAM[5982] = 8'b1110110;
DRAM[5983] = 8'b1110110;
DRAM[5984] = 8'b1110111;
DRAM[5985] = 8'b1110111;
DRAM[5986] = 8'b1110111;
DRAM[5987] = 8'b1110111;
DRAM[5988] = 8'b1110111;
DRAM[5989] = 8'b1110111;
DRAM[5990] = 8'b1110111;
DRAM[5991] = 8'b1110111;
DRAM[5992] = 8'b1110111;
DRAM[5993] = 8'b1110111;
DRAM[5994] = 8'b1110111;
DRAM[5995] = 8'b1110111;
DRAM[5996] = 8'b1110111;
DRAM[5997] = 8'b1110111;
DRAM[5998] = 8'b1110111;
DRAM[5999] = 8'b1110111;
DRAM[6000] = 8'b1110100;
DRAM[6001] = 8'b1110101;
DRAM[6002] = 8'b1110101;
DRAM[6003] = 8'b1110110;
DRAM[6004] = 8'b1110110;
DRAM[6005] = 8'b1110111;
DRAM[6006] = 8'b1111000;
DRAM[6007] = 8'b1111000;
DRAM[6008] = 8'b1110011;
DRAM[6009] = 8'b1111000;
DRAM[6010] = 8'b1111110;
DRAM[6011] = 8'b10000010;
DRAM[6012] = 8'b10000100;
DRAM[6013] = 8'b10001000;
DRAM[6014] = 8'b10001110;
DRAM[6015] = 8'b10010011;
DRAM[6016] = 8'b1111011;
DRAM[6017] = 8'b1111001;
DRAM[6018] = 8'b1111000;
DRAM[6019] = 8'b1111011;
DRAM[6020] = 8'b1111111;
DRAM[6021] = 8'b1111111;
DRAM[6022] = 8'b1111001;
DRAM[6023] = 8'b1110100;
DRAM[6024] = 8'b1110110;
DRAM[6025] = 8'b1111000;
DRAM[6026] = 8'b1111011;
DRAM[6027] = 8'b1111101;
DRAM[6028] = 8'b1111100;
DRAM[6029] = 8'b1111001;
DRAM[6030] = 8'b1110101;
DRAM[6031] = 8'b1110011;
DRAM[6032] = 8'b1111010;
DRAM[6033] = 8'b1110001;
DRAM[6034] = 8'b10001011;
DRAM[6035] = 8'b1111010;
DRAM[6036] = 8'b1111011;
DRAM[6037] = 8'b10011000;
DRAM[6038] = 8'b10011011;
DRAM[6039] = 8'b11000000;
DRAM[6040] = 8'b10010111;
DRAM[6041] = 8'b10010011;
DRAM[6042] = 8'b10001011;
DRAM[6043] = 8'b10000001;
DRAM[6044] = 8'b1111000;
DRAM[6045] = 8'b1110101;
DRAM[6046] = 8'b1111000;
DRAM[6047] = 8'b1111100;
DRAM[6048] = 8'b1111010;
DRAM[6049] = 8'b1110101;
DRAM[6050] = 8'b1110010;
DRAM[6051] = 8'b1110010;
DRAM[6052] = 8'b1110110;
DRAM[6053] = 8'b1110111;
DRAM[6054] = 8'b1110011;
DRAM[6055] = 8'b1101110;
DRAM[6056] = 8'b1110001;
DRAM[6057] = 8'b1110001;
DRAM[6058] = 8'b1110000;
DRAM[6059] = 8'b1101111;
DRAM[6060] = 8'b1101111;
DRAM[6061] = 8'b1101110;
DRAM[6062] = 8'b1101101;
DRAM[6063] = 8'b1101101;
DRAM[6064] = 8'b1101100;
DRAM[6065] = 8'b1101100;
DRAM[6066] = 8'b1101100;
DRAM[6067] = 8'b1101011;
DRAM[6068] = 8'b1101011;
DRAM[6069] = 8'b1101010;
DRAM[6070] = 8'b1101010;
DRAM[6071] = 8'b1101010;
DRAM[6072] = 8'b1101001;
DRAM[6073] = 8'b1101001;
DRAM[6074] = 8'b1101000;
DRAM[6075] = 8'b1100111;
DRAM[6076] = 8'b1100101;
DRAM[6077] = 8'b1100100;
DRAM[6078] = 8'b1100011;
DRAM[6079] = 8'b1100011;
DRAM[6080] = 8'b1100010;
DRAM[6081] = 8'b1100010;
DRAM[6082] = 8'b1100011;
DRAM[6083] = 8'b1100010;
DRAM[6084] = 8'b1100001;
DRAM[6085] = 8'b1100000;
DRAM[6086] = 8'b1011111;
DRAM[6087] = 8'b1011110;
DRAM[6088] = 8'b1011111;
DRAM[6089] = 8'b1011111;
DRAM[6090] = 8'b1011110;
DRAM[6091] = 8'b1011110;
DRAM[6092] = 8'b1011101;
DRAM[6093] = 8'b1011100;
DRAM[6094] = 8'b1011011;
DRAM[6095] = 8'b1011011;
DRAM[6096] = 8'b1011001;
DRAM[6097] = 8'b1011000;
DRAM[6098] = 8'b1010111;
DRAM[6099] = 8'b1010110;
DRAM[6100] = 8'b1010110;
DRAM[6101] = 8'b1010110;
DRAM[6102] = 8'b1010110;
DRAM[6103] = 8'b1010111;
DRAM[6104] = 8'b1010101;
DRAM[6105] = 8'b1010101;
DRAM[6106] = 8'b1010101;
DRAM[6107] = 8'b1010100;
DRAM[6108] = 8'b1010100;
DRAM[6109] = 8'b1010011;
DRAM[6110] = 8'b1010011;
DRAM[6111] = 8'b1010011;
DRAM[6112] = 8'b1010001;
DRAM[6113] = 8'b1010001;
DRAM[6114] = 8'b1010001;
DRAM[6115] = 8'b1010000;
DRAM[6116] = 8'b1010000;
DRAM[6117] = 8'b1010000;
DRAM[6118] = 8'b1001111;
DRAM[6119] = 8'b1001111;
DRAM[6120] = 8'b1001110;
DRAM[6121] = 8'b1001110;
DRAM[6122] = 8'b1001110;
DRAM[6123] = 8'b1001101;
DRAM[6124] = 8'b1001101;
DRAM[6125] = 8'b1001100;
DRAM[6126] = 8'b1001100;
DRAM[6127] = 8'b1001100;
DRAM[6128] = 8'b1001011;
DRAM[6129] = 8'b1001011;
DRAM[6130] = 8'b1001011;
DRAM[6131] = 8'b1001010;
DRAM[6132] = 8'b1001010;
DRAM[6133] = 8'b1001001;
DRAM[6134] = 8'b1001001;
DRAM[6135] = 8'b1001001;
DRAM[6136] = 8'b1001000;
DRAM[6137] = 8'b1001001;
DRAM[6138] = 8'b1001001;
DRAM[6139] = 8'b1001001;
DRAM[6140] = 8'b1001001;
DRAM[6141] = 8'b1001000;
DRAM[6142] = 8'b1000111;
DRAM[6143] = 8'b1000110;
DRAM[6144] = 8'b1100011;
DRAM[6145] = 8'b1100100;
DRAM[6146] = 8'b1100101;
DRAM[6147] = 8'b1100110;
DRAM[6148] = 8'b1100110;
DRAM[6149] = 8'b1100100;
DRAM[6150] = 8'b1100011;
DRAM[6151] = 8'b1100010;
DRAM[6152] = 8'b1100101;
DRAM[6153] = 8'b1100101;
DRAM[6154] = 8'b1100101;
DRAM[6155] = 8'b1100110;
DRAM[6156] = 8'b1100110;
DRAM[6157] = 8'b1100111;
DRAM[6158] = 8'b1100111;
DRAM[6159] = 8'b1100111;
DRAM[6160] = 8'b1101000;
DRAM[6161] = 8'b1101001;
DRAM[6162] = 8'b1101010;
DRAM[6163] = 8'b1101011;
DRAM[6164] = 8'b1101101;
DRAM[6165] = 8'b1101110;
DRAM[6166] = 8'b1101111;
DRAM[6167] = 8'b1110000;
DRAM[6168] = 8'b1110000;
DRAM[6169] = 8'b1101111;
DRAM[6170] = 8'b1101111;
DRAM[6171] = 8'b1101111;
DRAM[6172] = 8'b1101111;
DRAM[6173] = 8'b1101111;
DRAM[6174] = 8'b1101110;
DRAM[6175] = 8'b1101110;
DRAM[6176] = 8'b1110000;
DRAM[6177] = 8'b1110000;
DRAM[6178] = 8'b1110000;
DRAM[6179] = 8'b1110001;
DRAM[6180] = 8'b1110001;
DRAM[6181] = 8'b1110010;
DRAM[6182] = 8'b1110010;
DRAM[6183] = 8'b1110010;
DRAM[6184] = 8'b1110011;
DRAM[6185] = 8'b1110011;
DRAM[6186] = 8'b1110011;
DRAM[6187] = 8'b1110011;
DRAM[6188] = 8'b1110011;
DRAM[6189] = 8'b1110011;
DRAM[6190] = 8'b1110011;
DRAM[6191] = 8'b1110011;
DRAM[6192] = 8'b1110010;
DRAM[6193] = 8'b1110011;
DRAM[6194] = 8'b1110100;
DRAM[6195] = 8'b1110101;
DRAM[6196] = 8'b1110101;
DRAM[6197] = 8'b1110101;
DRAM[6198] = 8'b1110101;
DRAM[6199] = 8'b1110100;
DRAM[6200] = 8'b1110001;
DRAM[6201] = 8'b1110010;
DRAM[6202] = 8'b1110100;
DRAM[6203] = 8'b1110110;
DRAM[6204] = 8'b1111000;
DRAM[6205] = 8'b1111001;
DRAM[6206] = 8'b1111001;
DRAM[6207] = 8'b1111001;
DRAM[6208] = 8'b1111000;
DRAM[6209] = 8'b1111000;
DRAM[6210] = 8'b1111000;
DRAM[6211] = 8'b1111000;
DRAM[6212] = 8'b1111000;
DRAM[6213] = 8'b1111000;
DRAM[6214] = 8'b1111000;
DRAM[6215] = 8'b1111000;
DRAM[6216] = 8'b1111010;
DRAM[6217] = 8'b1111010;
DRAM[6218] = 8'b1111001;
DRAM[6219] = 8'b1110111;
DRAM[6220] = 8'b1110111;
DRAM[6221] = 8'b1110111;
DRAM[6222] = 8'b1110111;
DRAM[6223] = 8'b1110111;
DRAM[6224] = 8'b1110100;
DRAM[6225] = 8'b1110101;
DRAM[6226] = 8'b1110110;
DRAM[6227] = 8'b1110111;
DRAM[6228] = 8'b1111000;
DRAM[6229] = 8'b1111000;
DRAM[6230] = 8'b1111000;
DRAM[6231] = 8'b1111000;
DRAM[6232] = 8'b1111000;
DRAM[6233] = 8'b1111000;
DRAM[6234] = 8'b1111000;
DRAM[6235] = 8'b1111000;
DRAM[6236] = 8'b1111000;
DRAM[6237] = 8'b1111000;
DRAM[6238] = 8'b1111000;
DRAM[6239] = 8'b1111000;
DRAM[6240] = 8'b1111011;
DRAM[6241] = 8'b1110110;
DRAM[6242] = 8'b1110101;
DRAM[6243] = 8'b1111000;
DRAM[6244] = 8'b1111001;
DRAM[6245] = 8'b1110110;
DRAM[6246] = 8'b1110101;
DRAM[6247] = 8'b1110111;
DRAM[6248] = 8'b1110101;
DRAM[6249] = 8'b1111000;
DRAM[6250] = 8'b1110111;
DRAM[6251] = 8'b1110100;
DRAM[6252] = 8'b1110111;
DRAM[6253] = 8'b1111011;
DRAM[6254] = 8'b1111001;
DRAM[6255] = 8'b1110010;
DRAM[6256] = 8'b1110111;
DRAM[6257] = 8'b1111110;
DRAM[6258] = 8'b1110011;
DRAM[6259] = 8'b10000110;
DRAM[6260] = 8'b1110000;
DRAM[6261] = 8'b1101110;
DRAM[6262] = 8'b1110101;
DRAM[6263] = 8'b10001000;
DRAM[6264] = 8'b10000001;
DRAM[6265] = 8'b10000011;
DRAM[6266] = 8'b1110001;
DRAM[6267] = 8'b10101101;
DRAM[6268] = 8'b10101110;
DRAM[6269] = 8'b10110101;
DRAM[6270] = 8'b11001001;
DRAM[6271] = 8'b10111010;
DRAM[6272] = 8'b10100001;
DRAM[6273] = 8'b10100010;
DRAM[6274] = 8'b11001111;
DRAM[6275] = 8'b11011000;
DRAM[6276] = 8'b10100010;
DRAM[6277] = 8'b10011000;
DRAM[6278] = 8'b10101011;
DRAM[6279] = 8'b10011001;
DRAM[6280] = 8'b10110000;
DRAM[6281] = 8'b10001110;
DRAM[6282] = 8'b10011110;
DRAM[6283] = 8'b10001001;
DRAM[6284] = 8'b1110111;
DRAM[6285] = 8'b1111110;
DRAM[6286] = 8'b1110010;
DRAM[6287] = 8'b10001010;
DRAM[6288] = 8'b10010000;
DRAM[6289] = 8'b10010001;
DRAM[6290] = 8'b10101110;
DRAM[6291] = 8'b10111111;
DRAM[6292] = 8'b10111101;
DRAM[6293] = 8'b11010101;
DRAM[6294] = 8'b11100111;
DRAM[6295] = 8'b11010010;
DRAM[6296] = 8'b11011000;
DRAM[6297] = 8'b11010100;
DRAM[6298] = 8'b10100010;
DRAM[6299] = 8'b1100111;
DRAM[6300] = 8'b1111101;
DRAM[6301] = 8'b10100000;
DRAM[6302] = 8'b10001110;
DRAM[6303] = 8'b10001010;
DRAM[6304] = 8'b1110011;
DRAM[6305] = 8'b10010001;
DRAM[6306] = 8'b1111011;
DRAM[6307] = 8'b1110011;
DRAM[6308] = 8'b1110111;
DRAM[6309] = 8'b1101111;
DRAM[6310] = 8'b1111001;
DRAM[6311] = 8'b1110111;
DRAM[6312] = 8'b1101111;
DRAM[6313] = 8'b1101111;
DRAM[6314] = 8'b1111000;
DRAM[6315] = 8'b1101000;
DRAM[6316] = 8'b1110011;
DRAM[6317] = 8'b1101001;
DRAM[6318] = 8'b1110011;
DRAM[6319] = 8'b1101100;
DRAM[6320] = 8'b1100110;
DRAM[6321] = 8'b1101011;
DRAM[6322] = 8'b1101011;
DRAM[6323] = 8'b1100111;
DRAM[6324] = 8'b1101000;
DRAM[6325] = 8'b1101101;
DRAM[6326] = 8'b1101101;
DRAM[6327] = 8'b1101001;
DRAM[6328] = 8'b1100111;
DRAM[6329] = 8'b1101000;
DRAM[6330] = 8'b1101000;
DRAM[6331] = 8'b1101000;
DRAM[6332] = 8'b1101000;
DRAM[6333] = 8'b1100111;
DRAM[6334] = 8'b1100110;
DRAM[6335] = 8'b1100101;
DRAM[6336] = 8'b1100010;
DRAM[6337] = 8'b1100010;
DRAM[6338] = 8'b1100011;
DRAM[6339] = 8'b1100011;
DRAM[6340] = 8'b1100011;
DRAM[6341] = 8'b1100010;
DRAM[6342] = 8'b1100001;
DRAM[6343] = 8'b1100001;
DRAM[6344] = 8'b1011111;
DRAM[6345] = 8'b1011111;
DRAM[6346] = 8'b1011110;
DRAM[6347] = 8'b1011101;
DRAM[6348] = 8'b1011101;
DRAM[6349] = 8'b1011100;
DRAM[6350] = 8'b1011011;
DRAM[6351] = 8'b1011011;
DRAM[6352] = 8'b1011001;
DRAM[6353] = 8'b1011001;
DRAM[6354] = 8'b1011000;
DRAM[6355] = 8'b1011000;
DRAM[6356] = 8'b1011000;
DRAM[6357] = 8'b1011000;
DRAM[6358] = 8'b1010111;
DRAM[6359] = 8'b1010111;
DRAM[6360] = 8'b1010101;
DRAM[6361] = 8'b1010101;
DRAM[6362] = 8'b1010101;
DRAM[6363] = 8'b1010100;
DRAM[6364] = 8'b1010100;
DRAM[6365] = 8'b1010011;
DRAM[6366] = 8'b1010011;
DRAM[6367] = 8'b1010011;
DRAM[6368] = 8'b1010010;
DRAM[6369] = 8'b1010010;
DRAM[6370] = 8'b1010010;
DRAM[6371] = 8'b1010001;
DRAM[6372] = 8'b1010001;
DRAM[6373] = 8'b1010000;
DRAM[6374] = 8'b1010000;
DRAM[6375] = 8'b1010000;
DRAM[6376] = 8'b1001111;
DRAM[6377] = 8'b1001111;
DRAM[6378] = 8'b1001111;
DRAM[6379] = 8'b1001110;
DRAM[6380] = 8'b1001110;
DRAM[6381] = 8'b1001101;
DRAM[6382] = 8'b1001101;
DRAM[6383] = 8'b1001101;
DRAM[6384] = 8'b1001101;
DRAM[6385] = 8'b1001101;
DRAM[6386] = 8'b1001101;
DRAM[6387] = 8'b1001100;
DRAM[6388] = 8'b1001100;
DRAM[6389] = 8'b1001011;
DRAM[6390] = 8'b1001011;
DRAM[6391] = 8'b1001011;
DRAM[6392] = 8'b1001010;
DRAM[6393] = 8'b1001010;
DRAM[6394] = 8'b1001010;
DRAM[6395] = 8'b1001001;
DRAM[6396] = 8'b1001001;
DRAM[6397] = 8'b1001000;
DRAM[6398] = 8'b1001000;
DRAM[6399] = 8'b1001000;
DRAM[6400] = 8'b1100011;
DRAM[6401] = 8'b1100011;
DRAM[6402] = 8'b1100101;
DRAM[6403] = 8'b1100101;
DRAM[6404] = 8'b1100101;
DRAM[6405] = 8'b1100100;
DRAM[6406] = 8'b1100011;
DRAM[6407] = 8'b1100010;
DRAM[6408] = 8'b1100101;
DRAM[6409] = 8'b1100101;
DRAM[6410] = 8'b1100110;
DRAM[6411] = 8'b1100110;
DRAM[6412] = 8'b1100110;
DRAM[6413] = 8'b1100111;
DRAM[6414] = 8'b1100111;
DRAM[6415] = 8'b1100111;
DRAM[6416] = 8'b1101001;
DRAM[6417] = 8'b1101001;
DRAM[6418] = 8'b1101010;
DRAM[6419] = 8'b1101011;
DRAM[6420] = 8'b1101101;
DRAM[6421] = 8'b1101110;
DRAM[6422] = 8'b1101111;
DRAM[6423] = 8'b1101111;
DRAM[6424] = 8'b1101111;
DRAM[6425] = 8'b1101111;
DRAM[6426] = 8'b1101111;
DRAM[6427] = 8'b1101111;
DRAM[6428] = 8'b1101111;
DRAM[6429] = 8'b1101111;
DRAM[6430] = 8'b1101111;
DRAM[6431] = 8'b1110000;
DRAM[6432] = 8'b1110000;
DRAM[6433] = 8'b1110000;
DRAM[6434] = 8'b1110001;
DRAM[6435] = 8'b1110001;
DRAM[6436] = 8'b1110001;
DRAM[6437] = 8'b1110010;
DRAM[6438] = 8'b1110010;
DRAM[6439] = 8'b1110010;
DRAM[6440] = 8'b1110011;
DRAM[6441] = 8'b1110011;
DRAM[6442] = 8'b1110011;
DRAM[6443] = 8'b1110011;
DRAM[6444] = 8'b1110011;
DRAM[6445] = 8'b1110011;
DRAM[6446] = 8'b1110011;
DRAM[6447] = 8'b1110011;
DRAM[6448] = 8'b1110010;
DRAM[6449] = 8'b1110011;
DRAM[6450] = 8'b1110100;
DRAM[6451] = 8'b1110101;
DRAM[6452] = 8'b1110101;
DRAM[6453] = 8'b1110101;
DRAM[6454] = 8'b1110101;
DRAM[6455] = 8'b1110100;
DRAM[6456] = 8'b1110010;
DRAM[6457] = 8'b1110011;
DRAM[6458] = 8'b1110101;
DRAM[6459] = 8'b1110110;
DRAM[6460] = 8'b1111000;
DRAM[6461] = 8'b1111000;
DRAM[6462] = 8'b1111000;
DRAM[6463] = 8'b1111000;
DRAM[6464] = 8'b1111000;
DRAM[6465] = 8'b1111000;
DRAM[6466] = 8'b1111000;
DRAM[6467] = 8'b1111000;
DRAM[6468] = 8'b1111000;
DRAM[6469] = 8'b1111000;
DRAM[6470] = 8'b1111000;
DRAM[6471] = 8'b1111000;
DRAM[6472] = 8'b1111010;
DRAM[6473] = 8'b1111001;
DRAM[6474] = 8'b1111000;
DRAM[6475] = 8'b1110111;
DRAM[6476] = 8'b1110111;
DRAM[6477] = 8'b1110111;
DRAM[6478] = 8'b1111000;
DRAM[6479] = 8'b1111000;
DRAM[6480] = 8'b1110110;
DRAM[6481] = 8'b1110110;
DRAM[6482] = 8'b1110111;
DRAM[6483] = 8'b1111000;
DRAM[6484] = 8'b1111000;
DRAM[6485] = 8'b1111000;
DRAM[6486] = 8'b1110111;
DRAM[6487] = 8'b1110111;
DRAM[6488] = 8'b1111000;
DRAM[6489] = 8'b1111000;
DRAM[6490] = 8'b1111000;
DRAM[6491] = 8'b1111000;
DRAM[6492] = 8'b1111000;
DRAM[6493] = 8'b1111000;
DRAM[6494] = 8'b1111000;
DRAM[6495] = 8'b1111000;
DRAM[6496] = 8'b1110000;
DRAM[6497] = 8'b1110001;
DRAM[6498] = 8'b1110110;
DRAM[6499] = 8'b1111100;
DRAM[6500] = 8'b1111101;
DRAM[6501] = 8'b1111001;
DRAM[6502] = 8'b1111000;
DRAM[6503] = 8'b1111011;
DRAM[6504] = 8'b1111011;
DRAM[6505] = 8'b1111000;
DRAM[6506] = 8'b1111010;
DRAM[6507] = 8'b1111100;
DRAM[6508] = 8'b1110101;
DRAM[6509] = 8'b1101110;
DRAM[6510] = 8'b1110111;
DRAM[6511] = 8'b10001000;
DRAM[6512] = 8'b1111011;
DRAM[6513] = 8'b1111100;
DRAM[6514] = 8'b1111001;
DRAM[6515] = 8'b1111011;
DRAM[6516] = 8'b1111101;
DRAM[6517] = 8'b10001110;
DRAM[6518] = 8'b10001000;
DRAM[6519] = 8'b10000100;
DRAM[6520] = 8'b10001111;
DRAM[6521] = 8'b11000011;
DRAM[6522] = 8'b10101110;
DRAM[6523] = 8'b11000101;
DRAM[6524] = 8'b11010110;
DRAM[6525] = 8'b11101100;
DRAM[6526] = 8'b11110110;
DRAM[6527] = 8'b11100100;
DRAM[6528] = 8'b11101100;
DRAM[6529] = 8'b11100110;
DRAM[6530] = 8'b11111111;
DRAM[6531] = 8'b11111111;
DRAM[6532] = 8'b11100000;
DRAM[6533] = 8'b11011111;
DRAM[6534] = 8'b11110001;
DRAM[6535] = 8'b11100110;
DRAM[6536] = 8'b11100010;
DRAM[6537] = 8'b11000011;
DRAM[6538] = 8'b11010001;
DRAM[6539] = 8'b10111101;
DRAM[6540] = 8'b10101010;
DRAM[6541] = 8'b10101110;
DRAM[6542] = 8'b10100001;
DRAM[6543] = 8'b10110110;
DRAM[6544] = 8'b11010110;
DRAM[6545] = 8'b11010100;
DRAM[6546] = 8'b11101001;
DRAM[6547] = 8'b11110011;
DRAM[6548] = 8'b11101011;
DRAM[6549] = 8'b11111100;
DRAM[6550] = 8'b11111111;
DRAM[6551] = 8'b11110100;
DRAM[6552] = 8'b11110000;
DRAM[6553] = 8'b11100101;
DRAM[6554] = 8'b11001011;
DRAM[6555] = 8'b10110010;
DRAM[6556] = 8'b10111010;
DRAM[6557] = 8'b10110011;
DRAM[6558] = 8'b10011100;
DRAM[6559] = 8'b10110000;
DRAM[6560] = 8'b10010110;
DRAM[6561] = 8'b10011100;
DRAM[6562] = 8'b10000000;
DRAM[6563] = 8'b1111000;
DRAM[6564] = 8'b1110111;
DRAM[6565] = 8'b1101110;
DRAM[6566] = 8'b1110011;
DRAM[6567] = 8'b1101010;
DRAM[6568] = 8'b1110011;
DRAM[6569] = 8'b1100011;
DRAM[6570] = 8'b1100110;
DRAM[6571] = 8'b1110000;
DRAM[6572] = 8'b1111011;
DRAM[6573] = 8'b1101100;
DRAM[6574] = 8'b1101010;
DRAM[6575] = 8'b1101100;
DRAM[6576] = 8'b1101011;
DRAM[6577] = 8'b1101110;
DRAM[6578] = 8'b1101110;
DRAM[6579] = 8'b1101010;
DRAM[6580] = 8'b1101001;
DRAM[6581] = 8'b1101101;
DRAM[6582] = 8'b1101100;
DRAM[6583] = 8'b1101000;
DRAM[6584] = 8'b1100111;
DRAM[6585] = 8'b1101000;
DRAM[6586] = 8'b1101000;
DRAM[6587] = 8'b1101000;
DRAM[6588] = 8'b1101000;
DRAM[6589] = 8'b1100111;
DRAM[6590] = 8'b1100110;
DRAM[6591] = 8'b1100101;
DRAM[6592] = 8'b1100010;
DRAM[6593] = 8'b1100011;
DRAM[6594] = 8'b1100011;
DRAM[6595] = 8'b1100011;
DRAM[6596] = 8'b1100011;
DRAM[6597] = 8'b1100010;
DRAM[6598] = 8'b1100001;
DRAM[6599] = 8'b1100000;
DRAM[6600] = 8'b1011111;
DRAM[6601] = 8'b1011111;
DRAM[6602] = 8'b1011110;
DRAM[6603] = 8'b1011110;
DRAM[6604] = 8'b1011101;
DRAM[6605] = 8'b1011100;
DRAM[6606] = 8'b1011011;
DRAM[6607] = 8'b1011011;
DRAM[6608] = 8'b1011001;
DRAM[6609] = 8'b1011001;
DRAM[6610] = 8'b1011001;
DRAM[6611] = 8'b1011000;
DRAM[6612] = 8'b1011000;
DRAM[6613] = 8'b1011000;
DRAM[6614] = 8'b1010111;
DRAM[6615] = 8'b1010111;
DRAM[6616] = 8'b1010101;
DRAM[6617] = 8'b1010101;
DRAM[6618] = 8'b1010101;
DRAM[6619] = 8'b1010100;
DRAM[6620] = 8'b1010100;
DRAM[6621] = 8'b1010100;
DRAM[6622] = 8'b1010011;
DRAM[6623] = 8'b1010011;
DRAM[6624] = 8'b1010010;
DRAM[6625] = 8'b1010010;
DRAM[6626] = 8'b1010010;
DRAM[6627] = 8'b1010001;
DRAM[6628] = 8'b1010001;
DRAM[6629] = 8'b1010001;
DRAM[6630] = 8'b1010000;
DRAM[6631] = 8'b1010000;
DRAM[6632] = 8'b1001111;
DRAM[6633] = 8'b1001111;
DRAM[6634] = 8'b1001111;
DRAM[6635] = 8'b1001110;
DRAM[6636] = 8'b1001110;
DRAM[6637] = 8'b1001110;
DRAM[6638] = 8'b1001101;
DRAM[6639] = 8'b1001101;
DRAM[6640] = 8'b1001101;
DRAM[6641] = 8'b1001101;
DRAM[6642] = 8'b1001101;
DRAM[6643] = 8'b1001100;
DRAM[6644] = 8'b1001100;
DRAM[6645] = 8'b1001100;
DRAM[6646] = 8'b1001011;
DRAM[6647] = 8'b1001011;
DRAM[6648] = 8'b1001010;
DRAM[6649] = 8'b1001010;
DRAM[6650] = 8'b1001010;
DRAM[6651] = 8'b1001001;
DRAM[6652] = 8'b1001001;
DRAM[6653] = 8'b1001001;
DRAM[6654] = 8'b1001000;
DRAM[6655] = 8'b1001000;
DRAM[6656] = 8'b1100010;
DRAM[6657] = 8'b1100011;
DRAM[6658] = 8'b1100100;
DRAM[6659] = 8'b1100100;
DRAM[6660] = 8'b1100101;
DRAM[6661] = 8'b1100100;
DRAM[6662] = 8'b1100011;
DRAM[6663] = 8'b1100011;
DRAM[6664] = 8'b1100101;
DRAM[6665] = 8'b1100110;
DRAM[6666] = 8'b1100110;
DRAM[6667] = 8'b1100110;
DRAM[6668] = 8'b1100111;
DRAM[6669] = 8'b1100111;
DRAM[6670] = 8'b1100111;
DRAM[6671] = 8'b1100111;
DRAM[6672] = 8'b1101001;
DRAM[6673] = 8'b1101010;
DRAM[6674] = 8'b1101010;
DRAM[6675] = 8'b1101011;
DRAM[6676] = 8'b1101101;
DRAM[6677] = 8'b1101110;
DRAM[6678] = 8'b1101110;
DRAM[6679] = 8'b1101111;
DRAM[6680] = 8'b1101110;
DRAM[6681] = 8'b1101110;
DRAM[6682] = 8'b1101110;
DRAM[6683] = 8'b1101111;
DRAM[6684] = 8'b1110000;
DRAM[6685] = 8'b1110000;
DRAM[6686] = 8'b1110001;
DRAM[6687] = 8'b1110001;
DRAM[6688] = 8'b1110000;
DRAM[6689] = 8'b1110001;
DRAM[6690] = 8'b1110001;
DRAM[6691] = 8'b1110001;
DRAM[6692] = 8'b1110010;
DRAM[6693] = 8'b1110010;
DRAM[6694] = 8'b1110010;
DRAM[6695] = 8'b1110010;
DRAM[6696] = 8'b1110011;
DRAM[6697] = 8'b1110011;
DRAM[6698] = 8'b1110011;
DRAM[6699] = 8'b1110011;
DRAM[6700] = 8'b1110011;
DRAM[6701] = 8'b1110011;
DRAM[6702] = 8'b1110011;
DRAM[6703] = 8'b1110011;
DRAM[6704] = 8'b1110011;
DRAM[6705] = 8'b1110011;
DRAM[6706] = 8'b1110100;
DRAM[6707] = 8'b1110101;
DRAM[6708] = 8'b1110101;
DRAM[6709] = 8'b1110101;
DRAM[6710] = 8'b1110101;
DRAM[6711] = 8'b1110101;
DRAM[6712] = 8'b1110100;
DRAM[6713] = 8'b1110101;
DRAM[6714] = 8'b1110110;
DRAM[6715] = 8'b1110111;
DRAM[6716] = 8'b1110111;
DRAM[6717] = 8'b1110111;
DRAM[6718] = 8'b1110111;
DRAM[6719] = 8'b1110111;
DRAM[6720] = 8'b1111000;
DRAM[6721] = 8'b1111000;
DRAM[6722] = 8'b1111000;
DRAM[6723] = 8'b1111000;
DRAM[6724] = 8'b1111000;
DRAM[6725] = 8'b1111000;
DRAM[6726] = 8'b1111000;
DRAM[6727] = 8'b1111000;
DRAM[6728] = 8'b1111001;
DRAM[6729] = 8'b1111000;
DRAM[6730] = 8'b1111000;
DRAM[6731] = 8'b1110111;
DRAM[6732] = 8'b1111000;
DRAM[6733] = 8'b1111000;
DRAM[6734] = 8'b1111001;
DRAM[6735] = 8'b1111010;
DRAM[6736] = 8'b1111000;
DRAM[6737] = 8'b1111000;
DRAM[6738] = 8'b1111001;
DRAM[6739] = 8'b1111001;
DRAM[6740] = 8'b1111000;
DRAM[6741] = 8'b1111000;
DRAM[6742] = 8'b1110111;
DRAM[6743] = 8'b1110110;
DRAM[6744] = 8'b1111000;
DRAM[6745] = 8'b1111000;
DRAM[6746] = 8'b1111000;
DRAM[6747] = 8'b1111000;
DRAM[6748] = 8'b1111000;
DRAM[6749] = 8'b1111001;
DRAM[6750] = 8'b1111001;
DRAM[6751] = 8'b1111001;
DRAM[6752] = 8'b1110100;
DRAM[6753] = 8'b1110100;
DRAM[6754] = 8'b1111000;
DRAM[6755] = 8'b1111011;
DRAM[6756] = 8'b1111000;
DRAM[6757] = 8'b1110011;
DRAM[6758] = 8'b1110100;
DRAM[6759] = 8'b1111001;
DRAM[6760] = 8'b10000000;
DRAM[6761] = 8'b1110010;
DRAM[6762] = 8'b1101100;
DRAM[6763] = 8'b1110111;
DRAM[6764] = 8'b10000011;
DRAM[6765] = 8'b10000001;
DRAM[6766] = 8'b1111000;
DRAM[6767] = 8'b1110010;
DRAM[6768] = 8'b10000101;
DRAM[6769] = 8'b10010000;
DRAM[6770] = 8'b10110001;
DRAM[6771] = 8'b10100100;
DRAM[6772] = 8'b10111101;
DRAM[6773] = 8'b11011110;
DRAM[6774] = 8'b11010001;
DRAM[6775] = 8'b11000011;
DRAM[6776] = 8'b10110111;
DRAM[6777] = 8'b11111110;
DRAM[6778] = 8'b11100110;
DRAM[6779] = 8'b11100011;
DRAM[6780] = 8'b11111000;
DRAM[6781] = 8'b11111111;
DRAM[6782] = 8'b11111111;
DRAM[6783] = 8'b11111100;
DRAM[6784] = 8'b11111111;
DRAM[6785] = 8'b11111001;
DRAM[6786] = 8'b11111110;
DRAM[6787] = 8'b11111111;
DRAM[6788] = 8'b11110110;
DRAM[6789] = 8'b11111010;
DRAM[6790] = 8'b11111111;
DRAM[6791] = 8'b11111101;
DRAM[6792] = 8'b11111111;
DRAM[6793] = 8'b11101001;
DRAM[6794] = 8'b11111001;
DRAM[6795] = 8'b11101110;
DRAM[6796] = 8'b11100010;
DRAM[6797] = 8'b11101001;
DRAM[6798] = 8'b11100001;
DRAM[6799] = 8'b11110001;
DRAM[6800] = 8'b11110100;
DRAM[6801] = 8'b11110000;
DRAM[6802] = 8'b11111100;
DRAM[6803] = 8'b11111110;
DRAM[6804] = 8'b11110011;
DRAM[6805] = 8'b11111101;
DRAM[6806] = 8'b11111111;
DRAM[6807] = 8'b11110010;
DRAM[6808] = 8'b11111111;
DRAM[6809] = 8'b11111000;
DRAM[6810] = 8'b11110100;
DRAM[6811] = 8'b11110001;
DRAM[6812] = 8'b11110101;
DRAM[6813] = 8'b11011100;
DRAM[6814] = 8'b10111000;
DRAM[6815] = 8'b11001000;
DRAM[6816] = 8'b10100001;
DRAM[6817] = 8'b10010000;
DRAM[6818] = 8'b1111100;
DRAM[6819] = 8'b1111111;
DRAM[6820] = 8'b1111101;
DRAM[6821] = 8'b1111000;
DRAM[6822] = 8'b10000000;
DRAM[6823] = 8'b1110100;
DRAM[6824] = 8'b1110101;
DRAM[6825] = 8'b1110001;
DRAM[6826] = 8'b1101111;
DRAM[6827] = 8'b1111110;
DRAM[6828] = 8'b1111100;
DRAM[6829] = 8'b1111000;
DRAM[6830] = 8'b1101110;
DRAM[6831] = 8'b1110000;
DRAM[6832] = 8'b1101111;
DRAM[6833] = 8'b1110001;
DRAM[6834] = 8'b1110000;
DRAM[6835] = 8'b1101100;
DRAM[6836] = 8'b1101011;
DRAM[6837] = 8'b1101100;
DRAM[6838] = 8'b1101011;
DRAM[6839] = 8'b1101000;
DRAM[6840] = 8'b1101000;
DRAM[6841] = 8'b1101000;
DRAM[6842] = 8'b1101000;
DRAM[6843] = 8'b1101000;
DRAM[6844] = 8'b1101000;
DRAM[6845] = 8'b1100111;
DRAM[6846] = 8'b1100110;
DRAM[6847] = 8'b1100110;
DRAM[6848] = 8'b1100011;
DRAM[6849] = 8'b1100011;
DRAM[6850] = 8'b1100011;
DRAM[6851] = 8'b1100011;
DRAM[6852] = 8'b1100011;
DRAM[6853] = 8'b1100010;
DRAM[6854] = 8'b1100001;
DRAM[6855] = 8'b1100000;
DRAM[6856] = 8'b1011111;
DRAM[6857] = 8'b1011111;
DRAM[6858] = 8'b1011111;
DRAM[6859] = 8'b1011110;
DRAM[6860] = 8'b1011101;
DRAM[6861] = 8'b1011100;
DRAM[6862] = 8'b1011100;
DRAM[6863] = 8'b1011011;
DRAM[6864] = 8'b1011010;
DRAM[6865] = 8'b1011001;
DRAM[6866] = 8'b1011001;
DRAM[6867] = 8'b1011001;
DRAM[6868] = 8'b1011000;
DRAM[6869] = 8'b1011000;
DRAM[6870] = 8'b1010111;
DRAM[6871] = 8'b1010111;
DRAM[6872] = 8'b1010101;
DRAM[6873] = 8'b1010101;
DRAM[6874] = 8'b1010101;
DRAM[6875] = 8'b1010101;
DRAM[6876] = 8'b1010100;
DRAM[6877] = 8'b1010100;
DRAM[6878] = 8'b1010100;
DRAM[6879] = 8'b1010011;
DRAM[6880] = 8'b1010010;
DRAM[6881] = 8'b1010010;
DRAM[6882] = 8'b1010010;
DRAM[6883] = 8'b1010010;
DRAM[6884] = 8'b1010001;
DRAM[6885] = 8'b1010001;
DRAM[6886] = 8'b1010001;
DRAM[6887] = 8'b1010000;
DRAM[6888] = 8'b1001111;
DRAM[6889] = 8'b1001111;
DRAM[6890] = 8'b1001111;
DRAM[6891] = 8'b1001111;
DRAM[6892] = 8'b1001110;
DRAM[6893] = 8'b1001110;
DRAM[6894] = 8'b1001110;
DRAM[6895] = 8'b1001101;
DRAM[6896] = 8'b1001101;
DRAM[6897] = 8'b1001101;
DRAM[6898] = 8'b1001101;
DRAM[6899] = 8'b1001101;
DRAM[6900] = 8'b1001100;
DRAM[6901] = 8'b1001100;
DRAM[6902] = 8'b1001100;
DRAM[6903] = 8'b1001011;
DRAM[6904] = 8'b1001010;
DRAM[6905] = 8'b1001010;
DRAM[6906] = 8'b1001010;
DRAM[6907] = 8'b1001010;
DRAM[6908] = 8'b1001001;
DRAM[6909] = 8'b1001001;
DRAM[6910] = 8'b1001001;
DRAM[6911] = 8'b1001000;
DRAM[6912] = 8'b1100010;
DRAM[6913] = 8'b1100010;
DRAM[6914] = 8'b1100011;
DRAM[6915] = 8'b1100011;
DRAM[6916] = 8'b1100100;
DRAM[6917] = 8'b1100100;
DRAM[6918] = 8'b1100100;
DRAM[6919] = 8'b1100100;
DRAM[6920] = 8'b1100110;
DRAM[6921] = 8'b1100110;
DRAM[6922] = 8'b1100110;
DRAM[6923] = 8'b1100111;
DRAM[6924] = 8'b1100111;
DRAM[6925] = 8'b1100111;
DRAM[6926] = 8'b1101000;
DRAM[6927] = 8'b1101000;
DRAM[6928] = 8'b1101010;
DRAM[6929] = 8'b1101010;
DRAM[6930] = 8'b1101011;
DRAM[6931] = 8'b1101100;
DRAM[6932] = 8'b1101100;
DRAM[6933] = 8'b1101101;
DRAM[6934] = 8'b1101110;
DRAM[6935] = 8'b1101110;
DRAM[6936] = 8'b1101101;
DRAM[6937] = 8'b1101110;
DRAM[6938] = 8'b1101110;
DRAM[6939] = 8'b1101111;
DRAM[6940] = 8'b1110000;
DRAM[6941] = 8'b1110001;
DRAM[6942] = 8'b1110010;
DRAM[6943] = 8'b1110010;
DRAM[6944] = 8'b1110001;
DRAM[6945] = 8'b1110001;
DRAM[6946] = 8'b1110001;
DRAM[6947] = 8'b1110010;
DRAM[6948] = 8'b1110010;
DRAM[6949] = 8'b1110010;
DRAM[6950] = 8'b1110011;
DRAM[6951] = 8'b1110011;
DRAM[6952] = 8'b1110100;
DRAM[6953] = 8'b1110100;
DRAM[6954] = 8'b1110100;
DRAM[6955] = 8'b1110100;
DRAM[6956] = 8'b1110100;
DRAM[6957] = 8'b1110100;
DRAM[6958] = 8'b1110100;
DRAM[6959] = 8'b1110100;
DRAM[6960] = 8'b1110011;
DRAM[6961] = 8'b1110100;
DRAM[6962] = 8'b1110101;
DRAM[6963] = 8'b1110101;
DRAM[6964] = 8'b1110110;
DRAM[6965] = 8'b1110110;
DRAM[6966] = 8'b1110101;
DRAM[6967] = 8'b1110101;
DRAM[6968] = 8'b1110110;
DRAM[6969] = 8'b1110111;
DRAM[6970] = 8'b1110111;
DRAM[6971] = 8'b1111000;
DRAM[6972] = 8'b1111000;
DRAM[6973] = 8'b1110111;
DRAM[6974] = 8'b1110110;
DRAM[6975] = 8'b1110110;
DRAM[6976] = 8'b1111001;
DRAM[6977] = 8'b1111001;
DRAM[6978] = 8'b1111001;
DRAM[6979] = 8'b1111001;
DRAM[6980] = 8'b1111001;
DRAM[6981] = 8'b1111001;
DRAM[6982] = 8'b1111001;
DRAM[6983] = 8'b1111001;
DRAM[6984] = 8'b1111000;
DRAM[6985] = 8'b1111000;
DRAM[6986] = 8'b1111000;
DRAM[6987] = 8'b1111000;
DRAM[6988] = 8'b1111000;
DRAM[6989] = 8'b1111001;
DRAM[6990] = 8'b1111010;
DRAM[6991] = 8'b1111011;
DRAM[6992] = 8'b1111001;
DRAM[6993] = 8'b1111010;
DRAM[6994] = 8'b1111010;
DRAM[6995] = 8'b1111010;
DRAM[6996] = 8'b1111001;
DRAM[6997] = 8'b1111000;
DRAM[6998] = 8'b1110111;
DRAM[6999] = 8'b1110110;
DRAM[7000] = 8'b1111000;
DRAM[7001] = 8'b1111000;
DRAM[7002] = 8'b1111000;
DRAM[7003] = 8'b1111001;
DRAM[7004] = 8'b1111001;
DRAM[7005] = 8'b1111001;
DRAM[7006] = 8'b1111001;
DRAM[7007] = 8'b1111010;
DRAM[7008] = 8'b10000000;
DRAM[7009] = 8'b1111010;
DRAM[7010] = 8'b1110110;
DRAM[7011] = 8'b1110110;
DRAM[7012] = 8'b1110110;
DRAM[7013] = 8'b1110101;
DRAM[7014] = 8'b1111000;
DRAM[7015] = 8'b1111110;
DRAM[7016] = 8'b1101101;
DRAM[7017] = 8'b1111111;
DRAM[7018] = 8'b10001010;
DRAM[7019] = 8'b10000001;
DRAM[7020] = 8'b1110010;
DRAM[7021] = 8'b1110000;
DRAM[7022] = 8'b1111011;
DRAM[7023] = 8'b10000101;
DRAM[7024] = 8'b10001001;
DRAM[7025] = 8'b10100001;
DRAM[7026] = 8'b11100111;
DRAM[7027] = 8'b11010100;
DRAM[7028] = 8'b11101100;
DRAM[7029] = 8'b11111111;
DRAM[7030] = 8'b11111011;
DRAM[7031] = 8'b11111001;
DRAM[7032] = 8'b11100101;
DRAM[7033] = 8'b11111111;
DRAM[7034] = 8'b11110101;
DRAM[7035] = 8'b11111011;
DRAM[7036] = 8'b11111111;
DRAM[7037] = 8'b11110111;
DRAM[7038] = 8'b11110110;
DRAM[7039] = 8'b11111111;
DRAM[7040] = 8'b11111001;
DRAM[7041] = 8'b11111001;
DRAM[7042] = 8'b11110111;
DRAM[7043] = 8'b11111001;
DRAM[7044] = 8'b11111111;
DRAM[7045] = 8'b11111111;
DRAM[7046] = 8'b11111010;
DRAM[7047] = 8'b11111001;
DRAM[7048] = 8'b11111111;
DRAM[7049] = 8'b11110010;
DRAM[7050] = 8'b11111111;
DRAM[7051] = 8'b11111111;
DRAM[7052] = 8'b11111010;
DRAM[7053] = 8'b11111111;
DRAM[7054] = 8'b11111111;
DRAM[7055] = 8'b11111111;
DRAM[7056] = 8'b11111100;
DRAM[7057] = 8'b11111000;
DRAM[7058] = 8'b11111110;
DRAM[7059] = 8'b11111110;
DRAM[7060] = 8'b11110101;
DRAM[7061] = 8'b11111011;
DRAM[7062] = 8'b11111111;
DRAM[7063] = 8'b11110100;
DRAM[7064] = 8'b11111111;
DRAM[7065] = 8'b11111111;
DRAM[7066] = 8'b11111111;
DRAM[7067] = 8'b11110111;
DRAM[7068] = 8'b11111111;
DRAM[7069] = 8'b11111111;
DRAM[7070] = 8'b11011010;
DRAM[7071] = 8'b11001001;
DRAM[7072] = 8'b10101110;
DRAM[7073] = 8'b10010110;
DRAM[7074] = 8'b10010010;
DRAM[7075] = 8'b10011000;
DRAM[7076] = 8'b10001000;
DRAM[7077] = 8'b1111101;
DRAM[7078] = 8'b10000011;
DRAM[7079] = 8'b1111011;
DRAM[7080] = 8'b1101100;
DRAM[7081] = 8'b10000011;
DRAM[7082] = 8'b1111110;
DRAM[7083] = 8'b1111010;
DRAM[7084] = 8'b1100101;
DRAM[7085] = 8'b1111000;
DRAM[7086] = 8'b1101111;
DRAM[7087] = 8'b1101001;
DRAM[7088] = 8'b1110000;
DRAM[7089] = 8'b1110000;
DRAM[7090] = 8'b1101111;
DRAM[7091] = 8'b1101101;
DRAM[7092] = 8'b1101100;
DRAM[7093] = 8'b1101100;
DRAM[7094] = 8'b1101011;
DRAM[7095] = 8'b1101010;
DRAM[7096] = 8'b1101000;
DRAM[7097] = 8'b1101000;
DRAM[7098] = 8'b1101001;
DRAM[7099] = 8'b1101001;
DRAM[7100] = 8'b1101000;
DRAM[7101] = 8'b1101000;
DRAM[7102] = 8'b1100111;
DRAM[7103] = 8'b1100110;
DRAM[7104] = 8'b1100100;
DRAM[7105] = 8'b1100100;
DRAM[7106] = 8'b1100100;
DRAM[7107] = 8'b1100100;
DRAM[7108] = 8'b1100011;
DRAM[7109] = 8'b1100010;
DRAM[7110] = 8'b1100001;
DRAM[7111] = 8'b1100000;
DRAM[7112] = 8'b1100000;
DRAM[7113] = 8'b1100000;
DRAM[7114] = 8'b1011111;
DRAM[7115] = 8'b1011110;
DRAM[7116] = 8'b1011101;
DRAM[7117] = 8'b1011101;
DRAM[7118] = 8'b1011100;
DRAM[7119] = 8'b1011100;
DRAM[7120] = 8'b1011011;
DRAM[7121] = 8'b1011010;
DRAM[7122] = 8'b1011010;
DRAM[7123] = 8'b1011001;
DRAM[7124] = 8'b1011000;
DRAM[7125] = 8'b1011000;
DRAM[7126] = 8'b1010111;
DRAM[7127] = 8'b1010111;
DRAM[7128] = 8'b1010110;
DRAM[7129] = 8'b1010110;
DRAM[7130] = 8'b1010101;
DRAM[7131] = 8'b1010101;
DRAM[7132] = 8'b1010101;
DRAM[7133] = 8'b1010100;
DRAM[7134] = 8'b1010100;
DRAM[7135] = 8'b1010100;
DRAM[7136] = 8'b1010011;
DRAM[7137] = 8'b1010011;
DRAM[7138] = 8'b1010010;
DRAM[7139] = 8'b1010010;
DRAM[7140] = 8'b1010010;
DRAM[7141] = 8'b1010001;
DRAM[7142] = 8'b1010001;
DRAM[7143] = 8'b1010001;
DRAM[7144] = 8'b1010000;
DRAM[7145] = 8'b1010000;
DRAM[7146] = 8'b1001111;
DRAM[7147] = 8'b1001111;
DRAM[7148] = 8'b1001111;
DRAM[7149] = 8'b1001110;
DRAM[7150] = 8'b1001110;
DRAM[7151] = 8'b1001110;
DRAM[7152] = 8'b1001110;
DRAM[7153] = 8'b1001110;
DRAM[7154] = 8'b1001101;
DRAM[7155] = 8'b1001101;
DRAM[7156] = 8'b1001101;
DRAM[7157] = 8'b1001100;
DRAM[7158] = 8'b1001100;
DRAM[7159] = 8'b1001100;
DRAM[7160] = 8'b1001011;
DRAM[7161] = 8'b1001011;
DRAM[7162] = 8'b1001010;
DRAM[7163] = 8'b1001010;
DRAM[7164] = 8'b1001010;
DRAM[7165] = 8'b1001001;
DRAM[7166] = 8'b1001001;
DRAM[7167] = 8'b1001001;
DRAM[7168] = 8'b1100010;
DRAM[7169] = 8'b1100010;
DRAM[7170] = 8'b1100010;
DRAM[7171] = 8'b1100010;
DRAM[7172] = 8'b1100011;
DRAM[7173] = 8'b1100011;
DRAM[7174] = 8'b1100100;
DRAM[7175] = 8'b1100100;
DRAM[7176] = 8'b1100110;
DRAM[7177] = 8'b1100110;
DRAM[7178] = 8'b1100111;
DRAM[7179] = 8'b1100111;
DRAM[7180] = 8'b1100111;
DRAM[7181] = 8'b1101000;
DRAM[7182] = 8'b1101000;
DRAM[7183] = 8'b1101000;
DRAM[7184] = 8'b1101010;
DRAM[7185] = 8'b1101010;
DRAM[7186] = 8'b1101011;
DRAM[7187] = 8'b1101100;
DRAM[7188] = 8'b1101100;
DRAM[7189] = 8'b1101101;
DRAM[7190] = 8'b1101110;
DRAM[7191] = 8'b1101110;
DRAM[7192] = 8'b1101110;
DRAM[7193] = 8'b1101110;
DRAM[7194] = 8'b1101111;
DRAM[7195] = 8'b1110000;
DRAM[7196] = 8'b1110001;
DRAM[7197] = 8'b1110010;
DRAM[7198] = 8'b1110010;
DRAM[7199] = 8'b1110011;
DRAM[7200] = 8'b1110001;
DRAM[7201] = 8'b1110001;
DRAM[7202] = 8'b1110010;
DRAM[7203] = 8'b1110010;
DRAM[7204] = 8'b1110010;
DRAM[7205] = 8'b1110011;
DRAM[7206] = 8'b1110011;
DRAM[7207] = 8'b1110011;
DRAM[7208] = 8'b1110100;
DRAM[7209] = 8'b1110100;
DRAM[7210] = 8'b1110100;
DRAM[7211] = 8'b1110100;
DRAM[7212] = 8'b1110100;
DRAM[7213] = 8'b1110100;
DRAM[7214] = 8'b1110100;
DRAM[7215] = 8'b1110100;
DRAM[7216] = 8'b1110011;
DRAM[7217] = 8'b1110100;
DRAM[7218] = 8'b1110101;
DRAM[7219] = 8'b1110110;
DRAM[7220] = 8'b1110110;
DRAM[7221] = 8'b1110110;
DRAM[7222] = 8'b1110110;
DRAM[7223] = 8'b1110101;
DRAM[7224] = 8'b1110111;
DRAM[7225] = 8'b1111000;
DRAM[7226] = 8'b1111000;
DRAM[7227] = 8'b1111000;
DRAM[7228] = 8'b1111000;
DRAM[7229] = 8'b1110111;
DRAM[7230] = 8'b1110110;
DRAM[7231] = 8'b1110110;
DRAM[7232] = 8'b1111001;
DRAM[7233] = 8'b1111001;
DRAM[7234] = 8'b1111001;
DRAM[7235] = 8'b1111001;
DRAM[7236] = 8'b1111001;
DRAM[7237] = 8'b1111001;
DRAM[7238] = 8'b1111001;
DRAM[7239] = 8'b1111001;
DRAM[7240] = 8'b1111000;
DRAM[7241] = 8'b1111000;
DRAM[7242] = 8'b1111000;
DRAM[7243] = 8'b1111000;
DRAM[7244] = 8'b1111001;
DRAM[7245] = 8'b1111010;
DRAM[7246] = 8'b1111011;
DRAM[7247] = 8'b1111100;
DRAM[7248] = 8'b1111010;
DRAM[7249] = 8'b1111010;
DRAM[7250] = 8'b1111011;
DRAM[7251] = 8'b1111011;
DRAM[7252] = 8'b1111010;
DRAM[7253] = 8'b1111001;
DRAM[7254] = 8'b1111000;
DRAM[7255] = 8'b1110111;
DRAM[7256] = 8'b1111000;
DRAM[7257] = 8'b1111000;
DRAM[7258] = 8'b1111000;
DRAM[7259] = 8'b1111001;
DRAM[7260] = 8'b1111001;
DRAM[7261] = 8'b1111010;
DRAM[7262] = 8'b1111010;
DRAM[7263] = 8'b1111011;
DRAM[7264] = 8'b10000000;
DRAM[7265] = 8'b1111001;
DRAM[7266] = 8'b1110101;
DRAM[7267] = 8'b1111000;
DRAM[7268] = 8'b1111101;
DRAM[7269] = 8'b1111111;
DRAM[7270] = 8'b10000000;
DRAM[7271] = 8'b10000011;
DRAM[7272] = 8'b1110000;
DRAM[7273] = 8'b1110100;
DRAM[7274] = 8'b1111011;
DRAM[7275] = 8'b10000000;
DRAM[7276] = 8'b1111100;
DRAM[7277] = 8'b1111101;
DRAM[7278] = 8'b10010000;
DRAM[7279] = 8'b10100111;
DRAM[7280] = 8'b10110101;
DRAM[7281] = 8'b11000011;
DRAM[7282] = 8'b11111111;
DRAM[7283] = 8'b11101111;
DRAM[7284] = 8'b11111001;
DRAM[7285] = 8'b11111111;
DRAM[7286] = 8'b11110101;
DRAM[7287] = 8'b11111111;
DRAM[7288] = 8'b11111111;
DRAM[7289] = 8'b11110100;
DRAM[7290] = 8'b11110110;
DRAM[7291] = 8'b11111111;
DRAM[7292] = 8'b11111111;
DRAM[7293] = 8'b11110100;
DRAM[7294] = 8'b11111111;
DRAM[7295] = 8'b11111111;
DRAM[7296] = 8'b11111110;
DRAM[7297] = 8'b11111111;
DRAM[7298] = 8'b11111111;
DRAM[7299] = 8'b11111111;
DRAM[7300] = 8'b11111111;
DRAM[7301] = 8'b11111111;
DRAM[7302] = 8'b11111101;
DRAM[7303] = 8'b11111111;
DRAM[7304] = 8'b11111111;
DRAM[7305] = 8'b11111001;
DRAM[7306] = 8'b11111111;
DRAM[7307] = 8'b11111111;
DRAM[7308] = 8'b11111011;
DRAM[7309] = 8'b11111110;
DRAM[7310] = 8'b11111110;
DRAM[7311] = 8'b11111111;
DRAM[7312] = 8'b11111111;
DRAM[7313] = 8'b11111111;
DRAM[7314] = 8'b11111111;
DRAM[7315] = 8'b11111111;
DRAM[7316] = 8'b11111110;
DRAM[7317] = 8'b11111111;
DRAM[7318] = 8'b11111111;
DRAM[7319] = 8'b11111111;
DRAM[7320] = 8'b11111010;
DRAM[7321] = 8'b11111111;
DRAM[7322] = 8'b11111111;
DRAM[7323] = 8'b11101111;
DRAM[7324] = 8'b11111010;
DRAM[7325] = 8'b11111111;
DRAM[7326] = 8'b11110010;
DRAM[7327] = 8'b11011101;
DRAM[7328] = 8'b11011101;
DRAM[7329] = 8'b11001001;
DRAM[7330] = 8'b11001111;
DRAM[7331] = 8'b11001000;
DRAM[7332] = 8'b10011110;
DRAM[7333] = 8'b10000000;
DRAM[7334] = 8'b1111001;
DRAM[7335] = 8'b1111000;
DRAM[7336] = 8'b10000011;
DRAM[7337] = 8'b10001110;
DRAM[7338] = 8'b1111110;
DRAM[7339] = 8'b1111000;
DRAM[7340] = 8'b1101000;
DRAM[7341] = 8'b1111101;
DRAM[7342] = 8'b1110011;
DRAM[7343] = 8'b1101101;
DRAM[7344] = 8'b1101110;
DRAM[7345] = 8'b1101101;
DRAM[7346] = 8'b1101101;
DRAM[7347] = 8'b1101101;
DRAM[7348] = 8'b1101101;
DRAM[7349] = 8'b1101100;
DRAM[7350] = 8'b1101011;
DRAM[7351] = 8'b1101100;
DRAM[7352] = 8'b1101000;
DRAM[7353] = 8'b1101001;
DRAM[7354] = 8'b1101001;
DRAM[7355] = 8'b1101001;
DRAM[7356] = 8'b1101001;
DRAM[7357] = 8'b1101000;
DRAM[7358] = 8'b1100111;
DRAM[7359] = 8'b1100110;
DRAM[7360] = 8'b1100101;
DRAM[7361] = 8'b1100101;
DRAM[7362] = 8'b1100101;
DRAM[7363] = 8'b1100101;
DRAM[7364] = 8'b1100100;
DRAM[7365] = 8'b1100010;
DRAM[7366] = 8'b1100001;
DRAM[7367] = 8'b1100000;
DRAM[7368] = 8'b1100000;
DRAM[7369] = 8'b1100000;
DRAM[7370] = 8'b1011111;
DRAM[7371] = 8'b1011111;
DRAM[7372] = 8'b1011110;
DRAM[7373] = 8'b1011101;
DRAM[7374] = 8'b1011100;
DRAM[7375] = 8'b1011100;
DRAM[7376] = 8'b1011100;
DRAM[7377] = 8'b1011011;
DRAM[7378] = 8'b1011011;
DRAM[7379] = 8'b1011010;
DRAM[7380] = 8'b1011001;
DRAM[7381] = 8'b1011000;
DRAM[7382] = 8'b1010111;
DRAM[7383] = 8'b1010111;
DRAM[7384] = 8'b1010110;
DRAM[7385] = 8'b1010110;
DRAM[7386] = 8'b1010110;
DRAM[7387] = 8'b1010101;
DRAM[7388] = 8'b1010101;
DRAM[7389] = 8'b1010101;
DRAM[7390] = 8'b1010100;
DRAM[7391] = 8'b1010100;
DRAM[7392] = 8'b1010011;
DRAM[7393] = 8'b1010011;
DRAM[7394] = 8'b1010011;
DRAM[7395] = 8'b1010010;
DRAM[7396] = 8'b1010010;
DRAM[7397] = 8'b1010010;
DRAM[7398] = 8'b1010001;
DRAM[7399] = 8'b1010001;
DRAM[7400] = 8'b1010000;
DRAM[7401] = 8'b1010000;
DRAM[7402] = 8'b1010000;
DRAM[7403] = 8'b1001111;
DRAM[7404] = 8'b1001111;
DRAM[7405] = 8'b1001111;
DRAM[7406] = 8'b1001110;
DRAM[7407] = 8'b1001110;
DRAM[7408] = 8'b1001110;
DRAM[7409] = 8'b1001110;
DRAM[7410] = 8'b1001110;
DRAM[7411] = 8'b1001101;
DRAM[7412] = 8'b1001101;
DRAM[7413] = 8'b1001101;
DRAM[7414] = 8'b1001100;
DRAM[7415] = 8'b1001100;
DRAM[7416] = 8'b1001011;
DRAM[7417] = 8'b1001011;
DRAM[7418] = 8'b1001011;
DRAM[7419] = 8'b1001010;
DRAM[7420] = 8'b1001010;
DRAM[7421] = 8'b1001010;
DRAM[7422] = 8'b1001001;
DRAM[7423] = 8'b1001001;
DRAM[7424] = 8'b1100001;
DRAM[7425] = 8'b1100001;
DRAM[7426] = 8'b1100001;
DRAM[7427] = 8'b1100001;
DRAM[7428] = 8'b1100010;
DRAM[7429] = 8'b1100011;
DRAM[7430] = 8'b1100100;
DRAM[7431] = 8'b1100101;
DRAM[7432] = 8'b1100111;
DRAM[7433] = 8'b1100111;
DRAM[7434] = 8'b1100111;
DRAM[7435] = 8'b1100111;
DRAM[7436] = 8'b1101000;
DRAM[7437] = 8'b1101000;
DRAM[7438] = 8'b1101000;
DRAM[7439] = 8'b1101001;
DRAM[7440] = 8'b1101011;
DRAM[7441] = 8'b1101011;
DRAM[7442] = 8'b1101011;
DRAM[7443] = 8'b1101100;
DRAM[7444] = 8'b1101100;
DRAM[7445] = 8'b1101101;
DRAM[7446] = 8'b1101101;
DRAM[7447] = 8'b1101101;
DRAM[7448] = 8'b1101111;
DRAM[7449] = 8'b1101111;
DRAM[7450] = 8'b1110000;
DRAM[7451] = 8'b1110000;
DRAM[7452] = 8'b1110001;
DRAM[7453] = 8'b1110010;
DRAM[7454] = 8'b1110010;
DRAM[7455] = 8'b1110010;
DRAM[7456] = 8'b1110010;
DRAM[7457] = 8'b1110010;
DRAM[7458] = 8'b1110010;
DRAM[7459] = 8'b1110010;
DRAM[7460] = 8'b1110011;
DRAM[7461] = 8'b1110011;
DRAM[7462] = 8'b1110011;
DRAM[7463] = 8'b1110100;
DRAM[7464] = 8'b1110101;
DRAM[7465] = 8'b1110101;
DRAM[7466] = 8'b1110101;
DRAM[7467] = 8'b1110101;
DRAM[7468] = 8'b1110101;
DRAM[7469] = 8'b1110101;
DRAM[7470] = 8'b1110101;
DRAM[7471] = 8'b1110101;
DRAM[7472] = 8'b1110100;
DRAM[7473] = 8'b1110100;
DRAM[7474] = 8'b1110101;
DRAM[7475] = 8'b1110110;
DRAM[7476] = 8'b1110111;
DRAM[7477] = 8'b1110111;
DRAM[7478] = 8'b1110110;
DRAM[7479] = 8'b1110110;
DRAM[7480] = 8'b1110111;
DRAM[7481] = 8'b1111000;
DRAM[7482] = 8'b1111000;
DRAM[7483] = 8'b1111000;
DRAM[7484] = 8'b1111000;
DRAM[7485] = 8'b1111000;
DRAM[7486] = 8'b1110111;
DRAM[7487] = 8'b1110110;
DRAM[7488] = 8'b1111010;
DRAM[7489] = 8'b1111010;
DRAM[7490] = 8'b1111010;
DRAM[7491] = 8'b1111010;
DRAM[7492] = 8'b1111010;
DRAM[7493] = 8'b1111010;
DRAM[7494] = 8'b1111010;
DRAM[7495] = 8'b1111010;
DRAM[7496] = 8'b1111010;
DRAM[7497] = 8'b1111001;
DRAM[7498] = 8'b1111001;
DRAM[7499] = 8'b1111001;
DRAM[7500] = 8'b1111001;
DRAM[7501] = 8'b1111010;
DRAM[7502] = 8'b1111010;
DRAM[7503] = 8'b1111011;
DRAM[7504] = 8'b1111010;
DRAM[7505] = 8'b1111010;
DRAM[7506] = 8'b1111011;
DRAM[7507] = 8'b1111011;
DRAM[7508] = 8'b1111011;
DRAM[7509] = 8'b1111010;
DRAM[7510] = 8'b1111001;
DRAM[7511] = 8'b1111001;
DRAM[7512] = 8'b1111000;
DRAM[7513] = 8'b1111000;
DRAM[7514] = 8'b1111001;
DRAM[7515] = 8'b1111001;
DRAM[7516] = 8'b1111010;
DRAM[7517] = 8'b1111011;
DRAM[7518] = 8'b1111011;
DRAM[7519] = 8'b1111011;
DRAM[7520] = 8'b1111100;
DRAM[7521] = 8'b1111000;
DRAM[7522] = 8'b1110111;
DRAM[7523] = 8'b1111100;
DRAM[7524] = 8'b1111110;
DRAM[7525] = 8'b1111011;
DRAM[7526] = 8'b1111001;
DRAM[7527] = 8'b1111001;
DRAM[7528] = 8'b10011011;
DRAM[7529] = 8'b10000011;
DRAM[7530] = 8'b10001111;
DRAM[7531] = 8'b11000111;
DRAM[7532] = 8'b11101101;
DRAM[7533] = 8'b11101010;
DRAM[7534] = 8'b11100101;
DRAM[7535] = 8'b11110000;
DRAM[7536] = 8'b11110010;
DRAM[7537] = 8'b11101011;
DRAM[7538] = 8'b11111111;
DRAM[7539] = 8'b11111010;
DRAM[7540] = 8'b11111110;
DRAM[7541] = 8'b11111111;
DRAM[7542] = 8'b11110111;
DRAM[7543] = 8'b11111111;
DRAM[7544] = 8'b11111111;
DRAM[7545] = 8'b11110110;
DRAM[7546] = 8'b11111111;
DRAM[7547] = 8'b11111111;
DRAM[7548] = 8'b11111101;
DRAM[7549] = 8'b11111100;
DRAM[7550] = 8'b11111111;
DRAM[7551] = 8'b11111101;
DRAM[7552] = 8'b11111111;
DRAM[7553] = 8'b11111111;
DRAM[7554] = 8'b11111101;
DRAM[7555] = 8'b11111001;
DRAM[7556] = 8'b11111110;
DRAM[7557] = 8'b11111101;
DRAM[7558] = 8'b11111011;
DRAM[7559] = 8'b11111111;
DRAM[7560] = 8'b11111111;
DRAM[7561] = 8'b11111110;
DRAM[7562] = 8'b11111111;
DRAM[7563] = 8'b11111111;
DRAM[7564] = 8'b11111100;
DRAM[7565] = 8'b11111110;
DRAM[7566] = 8'b11111111;
DRAM[7567] = 8'b11111011;
DRAM[7568] = 8'b11111101;
DRAM[7569] = 8'b11111110;
DRAM[7570] = 8'b11111101;
DRAM[7571] = 8'b11111011;
DRAM[7572] = 8'b11111100;
DRAM[7573] = 8'b11111101;
DRAM[7574] = 8'b11111101;
DRAM[7575] = 8'b11111101;
DRAM[7576] = 8'b11111110;
DRAM[7577] = 8'b11111001;
DRAM[7578] = 8'b11111111;
DRAM[7579] = 8'b11111001;
DRAM[7580] = 8'b11110110;
DRAM[7581] = 8'b11111101;
DRAM[7582] = 8'b11111001;
DRAM[7583] = 8'b11111111;
DRAM[7584] = 8'b11111010;
DRAM[7585] = 8'b11110001;
DRAM[7586] = 8'b11111110;
DRAM[7587] = 8'b11101110;
DRAM[7588] = 8'b11000101;
DRAM[7589] = 8'b10100111;
DRAM[7590] = 8'b10010111;
DRAM[7591] = 8'b10100010;
DRAM[7592] = 8'b10101010;
DRAM[7593] = 8'b10001011;
DRAM[7594] = 8'b1101111;
DRAM[7595] = 8'b1111000;
DRAM[7596] = 8'b1111010;
DRAM[7597] = 8'b1111001;
DRAM[7598] = 8'b1101111;
DRAM[7599] = 8'b1110011;
DRAM[7600] = 8'b1101111;
DRAM[7601] = 8'b1101100;
DRAM[7602] = 8'b1101100;
DRAM[7603] = 8'b1101110;
DRAM[7604] = 8'b1101110;
DRAM[7605] = 8'b1101011;
DRAM[7606] = 8'b1101011;
DRAM[7607] = 8'b1101110;
DRAM[7608] = 8'b1101001;
DRAM[7609] = 8'b1101001;
DRAM[7610] = 8'b1101010;
DRAM[7611] = 8'b1101010;
DRAM[7612] = 8'b1101001;
DRAM[7613] = 8'b1101000;
DRAM[7614] = 8'b1100111;
DRAM[7615] = 8'b1100111;
DRAM[7616] = 8'b1100110;
DRAM[7617] = 8'b1100110;
DRAM[7618] = 8'b1100110;
DRAM[7619] = 8'b1100101;
DRAM[7620] = 8'b1100100;
DRAM[7621] = 8'b1100010;
DRAM[7622] = 8'b1100001;
DRAM[7623] = 8'b1100000;
DRAM[7624] = 8'b1100001;
DRAM[7625] = 8'b1100000;
DRAM[7626] = 8'b1100000;
DRAM[7627] = 8'b1011111;
DRAM[7628] = 8'b1011110;
DRAM[7629] = 8'b1011101;
DRAM[7630] = 8'b1011101;
DRAM[7631] = 8'b1011101;
DRAM[7632] = 8'b1011100;
DRAM[7633] = 8'b1011100;
DRAM[7634] = 8'b1011011;
DRAM[7635] = 8'b1011010;
DRAM[7636] = 8'b1011001;
DRAM[7637] = 8'b1011000;
DRAM[7638] = 8'b1010111;
DRAM[7639] = 8'b1010111;
DRAM[7640] = 8'b1010111;
DRAM[7641] = 8'b1010110;
DRAM[7642] = 8'b1010110;
DRAM[7643] = 8'b1010110;
DRAM[7644] = 8'b1010101;
DRAM[7645] = 8'b1010101;
DRAM[7646] = 8'b1010101;
DRAM[7647] = 8'b1010101;
DRAM[7648] = 8'b1010100;
DRAM[7649] = 8'b1010011;
DRAM[7650] = 8'b1010011;
DRAM[7651] = 8'b1010011;
DRAM[7652] = 8'b1010010;
DRAM[7653] = 8'b1010010;
DRAM[7654] = 8'b1010010;
DRAM[7655] = 8'b1010010;
DRAM[7656] = 8'b1010001;
DRAM[7657] = 8'b1010000;
DRAM[7658] = 8'b1010000;
DRAM[7659] = 8'b1010000;
DRAM[7660] = 8'b1001111;
DRAM[7661] = 8'b1001111;
DRAM[7662] = 8'b1001111;
DRAM[7663] = 8'b1001111;
DRAM[7664] = 8'b1001111;
DRAM[7665] = 8'b1001110;
DRAM[7666] = 8'b1001110;
DRAM[7667] = 8'b1001110;
DRAM[7668] = 8'b1001101;
DRAM[7669] = 8'b1001101;
DRAM[7670] = 8'b1001101;
DRAM[7671] = 8'b1001101;
DRAM[7672] = 8'b1001100;
DRAM[7673] = 8'b1001011;
DRAM[7674] = 8'b1001011;
DRAM[7675] = 8'b1001011;
DRAM[7676] = 8'b1001010;
DRAM[7677] = 8'b1001010;
DRAM[7678] = 8'b1001010;
DRAM[7679] = 8'b1001010;
DRAM[7680] = 8'b1100001;
DRAM[7681] = 8'b1100001;
DRAM[7682] = 8'b1100000;
DRAM[7683] = 8'b1100000;
DRAM[7684] = 8'b1100001;
DRAM[7685] = 8'b1100011;
DRAM[7686] = 8'b1100101;
DRAM[7687] = 8'b1100110;
DRAM[7688] = 8'b1100111;
DRAM[7689] = 8'b1100111;
DRAM[7690] = 8'b1100111;
DRAM[7691] = 8'b1101000;
DRAM[7692] = 8'b1101000;
DRAM[7693] = 8'b1101000;
DRAM[7694] = 8'b1101001;
DRAM[7695] = 8'b1101001;
DRAM[7696] = 8'b1101011;
DRAM[7697] = 8'b1101011;
DRAM[7698] = 8'b1101100;
DRAM[7699] = 8'b1101100;
DRAM[7700] = 8'b1101100;
DRAM[7701] = 8'b1101100;
DRAM[7702] = 8'b1101101;
DRAM[7703] = 8'b1101101;
DRAM[7704] = 8'b1110000;
DRAM[7705] = 8'b1110001;
DRAM[7706] = 8'b1110001;
DRAM[7707] = 8'b1110001;
DRAM[7708] = 8'b1110001;
DRAM[7709] = 8'b1110001;
DRAM[7710] = 8'b1110001;
DRAM[7711] = 8'b1110001;
DRAM[7712] = 8'b1110010;
DRAM[7713] = 8'b1110010;
DRAM[7714] = 8'b1110010;
DRAM[7715] = 8'b1110011;
DRAM[7716] = 8'b1110011;
DRAM[7717] = 8'b1110011;
DRAM[7718] = 8'b1110100;
DRAM[7719] = 8'b1110100;
DRAM[7720] = 8'b1110101;
DRAM[7721] = 8'b1110101;
DRAM[7722] = 8'b1110101;
DRAM[7723] = 8'b1110101;
DRAM[7724] = 8'b1110101;
DRAM[7725] = 8'b1110101;
DRAM[7726] = 8'b1110101;
DRAM[7727] = 8'b1110101;
DRAM[7728] = 8'b1110100;
DRAM[7729] = 8'b1110101;
DRAM[7730] = 8'b1110110;
DRAM[7731] = 8'b1110110;
DRAM[7732] = 8'b1110111;
DRAM[7733] = 8'b1110111;
DRAM[7734] = 8'b1110110;
DRAM[7735] = 8'b1110110;
DRAM[7736] = 8'b1110111;
DRAM[7737] = 8'b1110111;
DRAM[7738] = 8'b1111000;
DRAM[7739] = 8'b1111001;
DRAM[7740] = 8'b1111001;
DRAM[7741] = 8'b1111000;
DRAM[7742] = 8'b1111000;
DRAM[7743] = 8'b1111000;
DRAM[7744] = 8'b1111010;
DRAM[7745] = 8'b1111010;
DRAM[7746] = 8'b1111010;
DRAM[7747] = 8'b1111010;
DRAM[7748] = 8'b1111010;
DRAM[7749] = 8'b1111010;
DRAM[7750] = 8'b1111010;
DRAM[7751] = 8'b1111010;
DRAM[7752] = 8'b1111011;
DRAM[7753] = 8'b1111011;
DRAM[7754] = 8'b1111010;
DRAM[7755] = 8'b1111001;
DRAM[7756] = 8'b1111001;
DRAM[7757] = 8'b1111001;
DRAM[7758] = 8'b1111010;
DRAM[7759] = 8'b1111010;
DRAM[7760] = 8'b1111001;
DRAM[7761] = 8'b1111010;
DRAM[7762] = 8'b1111011;
DRAM[7763] = 8'b1111011;
DRAM[7764] = 8'b1111100;
DRAM[7765] = 8'b1111011;
DRAM[7766] = 8'b1111011;
DRAM[7767] = 8'b1111011;
DRAM[7768] = 8'b1111000;
DRAM[7769] = 8'b1111000;
DRAM[7770] = 8'b1111001;
DRAM[7771] = 8'b1111001;
DRAM[7772] = 8'b1111010;
DRAM[7773] = 8'b1111011;
DRAM[7774] = 8'b1111100;
DRAM[7775] = 8'b1111100;
DRAM[7776] = 8'b1111101;
DRAM[7777] = 8'b1111100;
DRAM[7778] = 8'b1111101;
DRAM[7779] = 8'b1111110;
DRAM[7780] = 8'b1111011;
DRAM[7781] = 8'b1111010;
DRAM[7782] = 8'b10000001;
DRAM[7783] = 8'b10001011;
DRAM[7784] = 8'b10001101;
DRAM[7785] = 8'b10100010;
DRAM[7786] = 8'b11001101;
DRAM[7787] = 8'b11110101;
DRAM[7788] = 8'b11111111;
DRAM[7789] = 8'b11110110;
DRAM[7790] = 8'b11110111;
DRAM[7791] = 8'b11111111;
DRAM[7792] = 8'b11111010;
DRAM[7793] = 8'b11111001;
DRAM[7794] = 8'b11110100;
DRAM[7795] = 8'b11110110;
DRAM[7796] = 8'b11110101;
DRAM[7797] = 8'b11111111;
DRAM[7798] = 8'b11111010;
DRAM[7799] = 8'b11111100;
DRAM[7800] = 8'b11111111;
DRAM[7801] = 8'b11111111;
DRAM[7802] = 8'b11111111;
DRAM[7803] = 8'b11110101;
DRAM[7804] = 8'b11111111;
DRAM[7805] = 8'b11111101;
DRAM[7806] = 8'b11111111;
DRAM[7807] = 8'b11111010;
DRAM[7808] = 8'b11111111;
DRAM[7809] = 8'b11111111;
DRAM[7810] = 8'b11111111;
DRAM[7811] = 8'b11111101;
DRAM[7812] = 8'b11111100;
DRAM[7813] = 8'b11111110;
DRAM[7814] = 8'b11111111;
DRAM[7815] = 8'b11111111;
DRAM[7816] = 8'b11111111;
DRAM[7817] = 8'b11111101;
DRAM[7818] = 8'b11111110;
DRAM[7819] = 8'b11111111;
DRAM[7820] = 8'b11111110;
DRAM[7821] = 8'b11111111;
DRAM[7822] = 8'b11111111;
DRAM[7823] = 8'b11111110;
DRAM[7824] = 8'b11111111;
DRAM[7825] = 8'b11111111;
DRAM[7826] = 8'b11111111;
DRAM[7827] = 8'b11111110;
DRAM[7828] = 8'b11111111;
DRAM[7829] = 8'b11111111;
DRAM[7830] = 8'b11111100;
DRAM[7831] = 8'b11111111;
DRAM[7832] = 8'b11111111;
DRAM[7833] = 8'b11110101;
DRAM[7834] = 8'b11111111;
DRAM[7835] = 8'b11111111;
DRAM[7836] = 8'b11111011;
DRAM[7837] = 8'b11111010;
DRAM[7838] = 8'b11111001;
DRAM[7839] = 8'b11111111;
DRAM[7840] = 8'b11110111;
DRAM[7841] = 8'b11110111;
DRAM[7842] = 8'b11111111;
DRAM[7843] = 8'b11110110;
DRAM[7844] = 8'b11101011;
DRAM[7845] = 8'b11100001;
DRAM[7846] = 8'b11010001;
DRAM[7847] = 8'b11100101;
DRAM[7848] = 8'b11000100;
DRAM[7849] = 8'b10011001;
DRAM[7850] = 8'b10000000;
DRAM[7851] = 8'b1111111;
DRAM[7852] = 8'b10000100;
DRAM[7853] = 8'b1101111;
DRAM[7854] = 8'b1101110;
DRAM[7855] = 8'b1110110;
DRAM[7856] = 8'b1110011;
DRAM[7857] = 8'b1101111;
DRAM[7858] = 8'b1101110;
DRAM[7859] = 8'b1110001;
DRAM[7860] = 8'b1110000;
DRAM[7861] = 8'b1101011;
DRAM[7862] = 8'b1101010;
DRAM[7863] = 8'b1101110;
DRAM[7864] = 8'b1101001;
DRAM[7865] = 8'b1101001;
DRAM[7866] = 8'b1101010;
DRAM[7867] = 8'b1101010;
DRAM[7868] = 8'b1101001;
DRAM[7869] = 8'b1101001;
DRAM[7870] = 8'b1101000;
DRAM[7871] = 8'b1100111;
DRAM[7872] = 8'b1100110;
DRAM[7873] = 8'b1100110;
DRAM[7874] = 8'b1100110;
DRAM[7875] = 8'b1100101;
DRAM[7876] = 8'b1100100;
DRAM[7877] = 8'b1100010;
DRAM[7878] = 8'b1100001;
DRAM[7879] = 8'b1100000;
DRAM[7880] = 8'b1100001;
DRAM[7881] = 8'b1100001;
DRAM[7882] = 8'b1100000;
DRAM[7883] = 8'b1011111;
DRAM[7884] = 8'b1011110;
DRAM[7885] = 8'b1011110;
DRAM[7886] = 8'b1011101;
DRAM[7887] = 8'b1011101;
DRAM[7888] = 8'b1011101;
DRAM[7889] = 8'b1011101;
DRAM[7890] = 8'b1011100;
DRAM[7891] = 8'b1011011;
DRAM[7892] = 8'b1011001;
DRAM[7893] = 8'b1011000;
DRAM[7894] = 8'b1010111;
DRAM[7895] = 8'b1010111;
DRAM[7896] = 8'b1010111;
DRAM[7897] = 8'b1010111;
DRAM[7898] = 8'b1010110;
DRAM[7899] = 8'b1010110;
DRAM[7900] = 8'b1010110;
DRAM[7901] = 8'b1010101;
DRAM[7902] = 8'b1010101;
DRAM[7903] = 8'b1010101;
DRAM[7904] = 8'b1010100;
DRAM[7905] = 8'b1010100;
DRAM[7906] = 8'b1010011;
DRAM[7907] = 8'b1010011;
DRAM[7908] = 8'b1010011;
DRAM[7909] = 8'b1010010;
DRAM[7910] = 8'b1010010;
DRAM[7911] = 8'b1010010;
DRAM[7912] = 8'b1010001;
DRAM[7913] = 8'b1010001;
DRAM[7914] = 8'b1010000;
DRAM[7915] = 8'b1010000;
DRAM[7916] = 8'b1010000;
DRAM[7917] = 8'b1001111;
DRAM[7918] = 8'b1001111;
DRAM[7919] = 8'b1001111;
DRAM[7920] = 8'b1001111;
DRAM[7921] = 8'b1001111;
DRAM[7922] = 8'b1001110;
DRAM[7923] = 8'b1001110;
DRAM[7924] = 8'b1001110;
DRAM[7925] = 8'b1001101;
DRAM[7926] = 8'b1001101;
DRAM[7927] = 8'b1001101;
DRAM[7928] = 8'b1001100;
DRAM[7929] = 8'b1001100;
DRAM[7930] = 8'b1001011;
DRAM[7931] = 8'b1001011;
DRAM[7932] = 8'b1001011;
DRAM[7933] = 8'b1001010;
DRAM[7934] = 8'b1001010;
DRAM[7935] = 8'b1001010;
DRAM[7936] = 8'b1100001;
DRAM[7937] = 8'b1100001;
DRAM[7938] = 8'b1100000;
DRAM[7939] = 8'b1100000;
DRAM[7940] = 8'b1100001;
DRAM[7941] = 8'b1100011;
DRAM[7942] = 8'b1100101;
DRAM[7943] = 8'b1100110;
DRAM[7944] = 8'b1100111;
DRAM[7945] = 8'b1100111;
DRAM[7946] = 8'b1100111;
DRAM[7947] = 8'b1101000;
DRAM[7948] = 8'b1101000;
DRAM[7949] = 8'b1101001;
DRAM[7950] = 8'b1101001;
DRAM[7951] = 8'b1101001;
DRAM[7952] = 8'b1101011;
DRAM[7953] = 8'b1101011;
DRAM[7954] = 8'b1101100;
DRAM[7955] = 8'b1101100;
DRAM[7956] = 8'b1101100;
DRAM[7957] = 8'b1101100;
DRAM[7958] = 8'b1101101;
DRAM[7959] = 8'b1101101;
DRAM[7960] = 8'b1110010;
DRAM[7961] = 8'b1110010;
DRAM[7962] = 8'b1110001;
DRAM[7963] = 8'b1110001;
DRAM[7964] = 8'b1110001;
DRAM[7965] = 8'b1110001;
DRAM[7966] = 8'b1110001;
DRAM[7967] = 8'b1110000;
DRAM[7968] = 8'b1110010;
DRAM[7969] = 8'b1110010;
DRAM[7970] = 8'b1110010;
DRAM[7971] = 8'b1110011;
DRAM[7972] = 8'b1110011;
DRAM[7973] = 8'b1110100;
DRAM[7974] = 8'b1110100;
DRAM[7975] = 8'b1110100;
DRAM[7976] = 8'b1110101;
DRAM[7977] = 8'b1110101;
DRAM[7978] = 8'b1110101;
DRAM[7979] = 8'b1110101;
DRAM[7980] = 8'b1110101;
DRAM[7981] = 8'b1110101;
DRAM[7982] = 8'b1110101;
DRAM[7983] = 8'b1110101;
DRAM[7984] = 8'b1110100;
DRAM[7985] = 8'b1110101;
DRAM[7986] = 8'b1110110;
DRAM[7987] = 8'b1110111;
DRAM[7988] = 8'b1110111;
DRAM[7989] = 8'b1110111;
DRAM[7990] = 8'b1110111;
DRAM[7991] = 8'b1110110;
DRAM[7992] = 8'b1110110;
DRAM[7993] = 8'b1110111;
DRAM[7994] = 8'b1111000;
DRAM[7995] = 8'b1111001;
DRAM[7996] = 8'b1111001;
DRAM[7997] = 8'b1111001;
DRAM[7998] = 8'b1111001;
DRAM[7999] = 8'b1111000;
DRAM[8000] = 8'b1111010;
DRAM[8001] = 8'b1111010;
DRAM[8002] = 8'b1111010;
DRAM[8003] = 8'b1111010;
DRAM[8004] = 8'b1111010;
DRAM[8005] = 8'b1111010;
DRAM[8006] = 8'b1111010;
DRAM[8007] = 8'b1111010;
DRAM[8008] = 8'b1111100;
DRAM[8009] = 8'b1111100;
DRAM[8010] = 8'b1111011;
DRAM[8011] = 8'b1111010;
DRAM[8012] = 8'b1111001;
DRAM[8013] = 8'b1111001;
DRAM[8014] = 8'b1111001;
DRAM[8015] = 8'b1111001;
DRAM[8016] = 8'b1111001;
DRAM[8017] = 8'b1111001;
DRAM[8018] = 8'b1111011;
DRAM[8019] = 8'b1111100;
DRAM[8020] = 8'b1111100;
DRAM[8021] = 8'b1111100;
DRAM[8022] = 8'b1111100;
DRAM[8023] = 8'b1111100;
DRAM[8024] = 8'b1111000;
DRAM[8025] = 8'b1111000;
DRAM[8026] = 8'b1111001;
DRAM[8027] = 8'b1111010;
DRAM[8028] = 8'b1111011;
DRAM[8029] = 8'b1111011;
DRAM[8030] = 8'b1111100;
DRAM[8031] = 8'b1111101;
DRAM[8032] = 8'b1111101;
DRAM[8033] = 8'b1111111;
DRAM[8034] = 8'b10000010;
DRAM[8035] = 8'b10000000;
DRAM[8036] = 8'b1111111;
DRAM[8037] = 8'b10001000;
DRAM[8038] = 8'b10100010;
DRAM[8039] = 8'b10111011;
DRAM[8040] = 8'b11000110;
DRAM[8041] = 8'b11101101;
DRAM[8042] = 8'b11111111;
DRAM[8043] = 8'b11110111;
DRAM[8044] = 8'b11110010;
DRAM[8045] = 8'b11111111;
DRAM[8046] = 8'b11111111;
DRAM[8047] = 8'b11110000;
DRAM[8048] = 8'b11110001;
DRAM[8049] = 8'b11111111;
DRAM[8050] = 8'b11110111;
DRAM[8051] = 8'b11111111;
DRAM[8052] = 8'b11110011;
DRAM[8053] = 8'b11111111;
DRAM[8054] = 8'b11111111;
DRAM[8055] = 8'b11111011;
DRAM[8056] = 8'b11110110;
DRAM[8057] = 8'b11111111;
DRAM[8058] = 8'b11111111;
DRAM[8059] = 8'b11110000;
DRAM[8060] = 8'b11111111;
DRAM[8061] = 8'b11111100;
DRAM[8062] = 8'b11110011;
DRAM[8063] = 8'b11111111;
DRAM[8064] = 8'b11111111;
DRAM[8065] = 8'b11111011;
DRAM[8066] = 8'b11111111;
DRAM[8067] = 8'b11111111;
DRAM[8068] = 8'b11111111;
DRAM[8069] = 8'b11111111;
DRAM[8070] = 8'b11111111;
DRAM[8071] = 8'b11111001;
DRAM[8072] = 8'b11111111;
DRAM[8073] = 8'b11111110;
DRAM[8074] = 8'b11111011;
DRAM[8075] = 8'b11111111;
DRAM[8076] = 8'b11111010;
DRAM[8077] = 8'b11111011;
DRAM[8078] = 8'b11111111;
DRAM[8079] = 8'b11110111;
DRAM[8080] = 8'b11111110;
DRAM[8081] = 8'b11111111;
DRAM[8082] = 8'b11111110;
DRAM[8083] = 8'b11111101;
DRAM[8084] = 8'b11111111;
DRAM[8085] = 8'b11111110;
DRAM[8086] = 8'b11111001;
DRAM[8087] = 8'b11111111;
DRAM[8088] = 8'b11111111;
DRAM[8089] = 8'b11110100;
DRAM[8090] = 8'b11111110;
DRAM[8091] = 8'b11111110;
DRAM[8092] = 8'b11111110;
DRAM[8093] = 8'b11111111;
DRAM[8094] = 8'b11111010;
DRAM[8095] = 8'b11110011;
DRAM[8096] = 8'b11111000;
DRAM[8097] = 8'b11111001;
DRAM[8098] = 8'b11111111;
DRAM[8099] = 8'b11110001;
DRAM[8100] = 8'b11111011;
DRAM[8101] = 8'b11111111;
DRAM[8102] = 8'b11101110;
DRAM[8103] = 8'b11111111;
DRAM[8104] = 8'b11101001;
DRAM[8105] = 8'b11010010;
DRAM[8106] = 8'b11000101;
DRAM[8107] = 8'b10100101;
DRAM[8108] = 8'b10011110;
DRAM[8109] = 8'b10000101;
DRAM[8110] = 8'b10010000;
DRAM[8111] = 8'b10010110;
DRAM[8112] = 8'b1111000;
DRAM[8113] = 8'b1110010;
DRAM[8114] = 8'b1110001;
DRAM[8115] = 8'b1110011;
DRAM[8116] = 8'b1110001;
DRAM[8117] = 8'b1101011;
DRAM[8118] = 8'b1101001;
DRAM[8119] = 8'b1101101;
DRAM[8120] = 8'b1101001;
DRAM[8121] = 8'b1101010;
DRAM[8122] = 8'b1101010;
DRAM[8123] = 8'b1101010;
DRAM[8124] = 8'b1101010;
DRAM[8125] = 8'b1101001;
DRAM[8126] = 8'b1101000;
DRAM[8127] = 8'b1100111;
DRAM[8128] = 8'b1100111;
DRAM[8129] = 8'b1100111;
DRAM[8130] = 8'b1100110;
DRAM[8131] = 8'b1100110;
DRAM[8132] = 8'b1100100;
DRAM[8133] = 8'b1100010;
DRAM[8134] = 8'b1100001;
DRAM[8135] = 8'b1100000;
DRAM[8136] = 8'b1100001;
DRAM[8137] = 8'b1100001;
DRAM[8138] = 8'b1100000;
DRAM[8139] = 8'b1011111;
DRAM[8140] = 8'b1011111;
DRAM[8141] = 8'b1011110;
DRAM[8142] = 8'b1011101;
DRAM[8143] = 8'b1011101;
DRAM[8144] = 8'b1011110;
DRAM[8145] = 8'b1011101;
DRAM[8146] = 8'b1011100;
DRAM[8147] = 8'b1011011;
DRAM[8148] = 8'b1011001;
DRAM[8149] = 8'b1011000;
DRAM[8150] = 8'b1010111;
DRAM[8151] = 8'b1010111;
DRAM[8152] = 8'b1010111;
DRAM[8153] = 8'b1010111;
DRAM[8154] = 8'b1010111;
DRAM[8155] = 8'b1010110;
DRAM[8156] = 8'b1010110;
DRAM[8157] = 8'b1010101;
DRAM[8158] = 8'b1010101;
DRAM[8159] = 8'b1010101;
DRAM[8160] = 8'b1010100;
DRAM[8161] = 8'b1010100;
DRAM[8162] = 8'b1010100;
DRAM[8163] = 8'b1010011;
DRAM[8164] = 8'b1010011;
DRAM[8165] = 8'b1010010;
DRAM[8166] = 8'b1010010;
DRAM[8167] = 8'b1010010;
DRAM[8168] = 8'b1010001;
DRAM[8169] = 8'b1010001;
DRAM[8170] = 8'b1010001;
DRAM[8171] = 8'b1010000;
DRAM[8172] = 8'b1010000;
DRAM[8173] = 8'b1001111;
DRAM[8174] = 8'b1001111;
DRAM[8175] = 8'b1001111;
DRAM[8176] = 8'b1001111;
DRAM[8177] = 8'b1001111;
DRAM[8178] = 8'b1001111;
DRAM[8179] = 8'b1001110;
DRAM[8180] = 8'b1001110;
DRAM[8181] = 8'b1001101;
DRAM[8182] = 8'b1001101;
DRAM[8183] = 8'b1001101;
DRAM[8184] = 8'b1001100;
DRAM[8185] = 8'b1001100;
DRAM[8186] = 8'b1001100;
DRAM[8187] = 8'b1001011;
DRAM[8188] = 8'b1001011;
DRAM[8189] = 8'b1001010;
DRAM[8190] = 8'b1001010;
DRAM[8191] = 8'b1001010;
DRAM[8192] = 8'b1100001;
DRAM[8193] = 8'b1100010;
DRAM[8194] = 8'b1100011;
DRAM[8195] = 8'b1100101;
DRAM[8196] = 8'b1100111;
DRAM[8197] = 8'b1100111;
DRAM[8198] = 8'b1101000;
DRAM[8199] = 8'b1101000;
DRAM[8200] = 8'b1101000;
DRAM[8201] = 8'b1101000;
DRAM[8202] = 8'b1101000;
DRAM[8203] = 8'b1101001;
DRAM[8204] = 8'b1101001;
DRAM[8205] = 8'b1101010;
DRAM[8206] = 8'b1101010;
DRAM[8207] = 8'b1101010;
DRAM[8208] = 8'b1101011;
DRAM[8209] = 8'b1101011;
DRAM[8210] = 8'b1101100;
DRAM[8211] = 8'b1101101;
DRAM[8212] = 8'b1101101;
DRAM[8213] = 8'b1101110;
DRAM[8214] = 8'b1101111;
DRAM[8215] = 8'b1101111;
DRAM[8216] = 8'b1110001;
DRAM[8217] = 8'b1110001;
DRAM[8218] = 8'b1110001;
DRAM[8219] = 8'b1110010;
DRAM[8220] = 8'b1110010;
DRAM[8221] = 8'b1110011;
DRAM[8222] = 8'b1110011;
DRAM[8223] = 8'b1110011;
DRAM[8224] = 8'b1110010;
DRAM[8225] = 8'b1110010;
DRAM[8226] = 8'b1110010;
DRAM[8227] = 8'b1110011;
DRAM[8228] = 8'b1110011;
DRAM[8229] = 8'b1110100;
DRAM[8230] = 8'b1110100;
DRAM[8231] = 8'b1110100;
DRAM[8232] = 8'b1110110;
DRAM[8233] = 8'b1110110;
DRAM[8234] = 8'b1110111;
DRAM[8235] = 8'b1110111;
DRAM[8236] = 8'b1110111;
DRAM[8237] = 8'b1110110;
DRAM[8238] = 8'b1110101;
DRAM[8239] = 8'b1110101;
DRAM[8240] = 8'b1110101;
DRAM[8241] = 8'b1110110;
DRAM[8242] = 8'b1110111;
DRAM[8243] = 8'b1111000;
DRAM[8244] = 8'b1111000;
DRAM[8245] = 8'b1111000;
DRAM[8246] = 8'b1110111;
DRAM[8247] = 8'b1110111;
DRAM[8248] = 8'b1111000;
DRAM[8249] = 8'b1111001;
DRAM[8250] = 8'b1111001;
DRAM[8251] = 8'b1111010;
DRAM[8252] = 8'b1111010;
DRAM[8253] = 8'b1111001;
DRAM[8254] = 8'b1111001;
DRAM[8255] = 8'b1111000;
DRAM[8256] = 8'b1111010;
DRAM[8257] = 8'b1111010;
DRAM[8258] = 8'b1111010;
DRAM[8259] = 8'b1111010;
DRAM[8260] = 8'b1111010;
DRAM[8261] = 8'b1111010;
DRAM[8262] = 8'b1111010;
DRAM[8263] = 8'b1111010;
DRAM[8264] = 8'b1111101;
DRAM[8265] = 8'b1111100;
DRAM[8266] = 8'b1111100;
DRAM[8267] = 8'b1111011;
DRAM[8268] = 8'b1111011;
DRAM[8269] = 8'b1111010;
DRAM[8270] = 8'b1111010;
DRAM[8271] = 8'b1111010;
DRAM[8272] = 8'b1111011;
DRAM[8273] = 8'b1111010;
DRAM[8274] = 8'b1111001;
DRAM[8275] = 8'b1111001;
DRAM[8276] = 8'b1111010;
DRAM[8277] = 8'b1111011;
DRAM[8278] = 8'b1111010;
DRAM[8279] = 8'b1111001;
DRAM[8280] = 8'b1110011;
DRAM[8281] = 8'b10000100;
DRAM[8282] = 8'b1101100;
DRAM[8283] = 8'b1110110;
DRAM[8284] = 8'b10001010;
DRAM[8285] = 8'b10011000;
DRAM[8286] = 8'b1110101;
DRAM[8287] = 8'b1110010;
DRAM[8288] = 8'b1111010;
DRAM[8289] = 8'b10000011;
DRAM[8290] = 8'b10010100;
DRAM[8291] = 8'b10101011;
DRAM[8292] = 8'b11000100;
DRAM[8293] = 8'b11011100;
DRAM[8294] = 8'b11101110;
DRAM[8295] = 8'b11110111;
DRAM[8296] = 8'b11111001;
DRAM[8297] = 8'b11111001;
DRAM[8298] = 8'b11111001;
DRAM[8299] = 8'b11111001;
DRAM[8300] = 8'b11111001;
DRAM[8301] = 8'b11111001;
DRAM[8302] = 8'b11111001;
DRAM[8303] = 8'b11111001;
DRAM[8304] = 8'b11111000;
DRAM[8305] = 8'b11111001;
DRAM[8306] = 8'b11111001;
DRAM[8307] = 8'b11111010;
DRAM[8308] = 8'b11111011;
DRAM[8309] = 8'b11111100;
DRAM[8310] = 8'b11111101;
DRAM[8311] = 8'b11111101;
DRAM[8312] = 8'b11111110;
DRAM[8313] = 8'b11111110;
DRAM[8314] = 8'b11111110;
DRAM[8315] = 8'b11111111;
DRAM[8316] = 8'b11111111;
DRAM[8317] = 8'b11111111;
DRAM[8318] = 8'b11111111;
DRAM[8319] = 8'b11111111;
DRAM[8320] = 8'b11111111;
DRAM[8321] = 8'b11111111;
DRAM[8322] = 8'b11111111;
DRAM[8323] = 8'b11111111;
DRAM[8324] = 8'b11111111;
DRAM[8325] = 8'b11111111;
DRAM[8326] = 8'b11111111;
DRAM[8327] = 8'b11111111;
DRAM[8328] = 8'b11111111;
DRAM[8329] = 8'b11111111;
DRAM[8330] = 8'b11111111;
DRAM[8331] = 8'b11111111;
DRAM[8332] = 8'b11111111;
DRAM[8333] = 8'b11111111;
DRAM[8334] = 8'b11111111;
DRAM[8335] = 8'b11111111;
DRAM[8336] = 8'b11111111;
DRAM[8337] = 8'b11111111;
DRAM[8338] = 8'b11111111;
DRAM[8339] = 8'b11111111;
DRAM[8340] = 8'b11111111;
DRAM[8341] = 8'b11111111;
DRAM[8342] = 8'b11111111;
DRAM[8343] = 8'b11111111;
DRAM[8344] = 8'b11111100;
DRAM[8345] = 8'b11111100;
DRAM[8346] = 8'b11111100;
DRAM[8347] = 8'b11111101;
DRAM[8348] = 8'b11111101;
DRAM[8349] = 8'b11111110;
DRAM[8350] = 8'b11111110;
DRAM[8351] = 8'b11111110;
DRAM[8352] = 8'b11111010;
DRAM[8353] = 8'b11111010;
DRAM[8354] = 8'b11111010;
DRAM[8355] = 8'b11111010;
DRAM[8356] = 8'b11111010;
DRAM[8357] = 8'b11111010;
DRAM[8358] = 8'b11111010;
DRAM[8359] = 8'b11111010;
DRAM[8360] = 8'b11111111;
DRAM[8361] = 8'b11110101;
DRAM[8362] = 8'b11100111;
DRAM[8363] = 8'b11100001;
DRAM[8364] = 8'b11100010;
DRAM[8365] = 8'b11010100;
DRAM[8366] = 8'b10110000;
DRAM[8367] = 8'b10001011;
DRAM[8368] = 8'b1111010;
DRAM[8369] = 8'b1111110;
DRAM[8370] = 8'b10010010;
DRAM[8371] = 8'b1110111;
DRAM[8372] = 8'b1110000;
DRAM[8373] = 8'b10000000;
DRAM[8374] = 8'b1101100;
DRAM[8375] = 8'b1101101;
DRAM[8376] = 8'b1110110;
DRAM[8377] = 8'b1101011;
DRAM[8378] = 8'b1100111;
DRAM[8379] = 8'b1101110;
DRAM[8380] = 8'b1110010;
DRAM[8381] = 8'b1101100;
DRAM[8382] = 8'b1100110;
DRAM[8383] = 8'b1100101;
DRAM[8384] = 8'b1101101;
DRAM[8385] = 8'b1100101;
DRAM[8386] = 8'b1100101;
DRAM[8387] = 8'b1100100;
DRAM[8388] = 8'b1011110;
DRAM[8389] = 8'b1100011;
DRAM[8390] = 8'b1101000;
DRAM[8391] = 8'b1100010;
DRAM[8392] = 8'b1100100;
DRAM[8393] = 8'b1100001;
DRAM[8394] = 8'b1011110;
DRAM[8395] = 8'b1011101;
DRAM[8396] = 8'b1011110;
DRAM[8397] = 8'b1011110;
DRAM[8398] = 8'b1011110;
DRAM[8399] = 8'b1011101;
DRAM[8400] = 8'b1011101;
DRAM[8401] = 8'b1011101;
DRAM[8402] = 8'b1011100;
DRAM[8403] = 8'b1011011;
DRAM[8404] = 8'b1011011;
DRAM[8405] = 8'b1011010;
DRAM[8406] = 8'b1011001;
DRAM[8407] = 8'b1011001;
DRAM[8408] = 8'b1011001;
DRAM[8409] = 8'b1011001;
DRAM[8410] = 8'b1011000;
DRAM[8411] = 8'b1010111;
DRAM[8412] = 8'b1010111;
DRAM[8413] = 8'b1010110;
DRAM[8414] = 8'b1010101;
DRAM[8415] = 8'b1010101;
DRAM[8416] = 8'b1010100;
DRAM[8417] = 8'b1010100;
DRAM[8418] = 8'b1010100;
DRAM[8419] = 8'b1010100;
DRAM[8420] = 8'b1010100;
DRAM[8421] = 8'b1010100;
DRAM[8422] = 8'b1010100;
DRAM[8423] = 8'b1010100;
DRAM[8424] = 8'b1010001;
DRAM[8425] = 8'b1010010;
DRAM[8426] = 8'b1010010;
DRAM[8427] = 8'b1010011;
DRAM[8428] = 8'b1010011;
DRAM[8429] = 8'b1010010;
DRAM[8430] = 8'b1010010;
DRAM[8431] = 8'b1010001;
DRAM[8432] = 8'b1001111;
DRAM[8433] = 8'b1001111;
DRAM[8434] = 8'b1001111;
DRAM[8435] = 8'b1001110;
DRAM[8436] = 8'b1001110;
DRAM[8437] = 8'b1001101;
DRAM[8438] = 8'b1001101;
DRAM[8439] = 8'b1001101;
DRAM[8440] = 8'b1001101;
DRAM[8441] = 8'b1001101;
DRAM[8442] = 8'b1001101;
DRAM[8443] = 8'b1001100;
DRAM[8444] = 8'b1001100;
DRAM[8445] = 8'b1001011;
DRAM[8446] = 8'b1001011;
DRAM[8447] = 8'b1001011;
DRAM[8448] = 8'b1100001;
DRAM[8449] = 8'b1100010;
DRAM[8450] = 8'b1100011;
DRAM[8451] = 8'b1100101;
DRAM[8452] = 8'b1100110;
DRAM[8453] = 8'b1100111;
DRAM[8454] = 8'b1100111;
DRAM[8455] = 8'b1100111;
DRAM[8456] = 8'b1101000;
DRAM[8457] = 8'b1101000;
DRAM[8458] = 8'b1101000;
DRAM[8459] = 8'b1101001;
DRAM[8460] = 8'b1101001;
DRAM[8461] = 8'b1101010;
DRAM[8462] = 8'b1101010;
DRAM[8463] = 8'b1101010;
DRAM[8464] = 8'b1101011;
DRAM[8465] = 8'b1101011;
DRAM[8466] = 8'b1101100;
DRAM[8467] = 8'b1101101;
DRAM[8468] = 8'b1101101;
DRAM[8469] = 8'b1101110;
DRAM[8470] = 8'b1101111;
DRAM[8471] = 8'b1101111;
DRAM[8472] = 8'b1110001;
DRAM[8473] = 8'b1110001;
DRAM[8474] = 8'b1110001;
DRAM[8475] = 8'b1110010;
DRAM[8476] = 8'b1110010;
DRAM[8477] = 8'b1110010;
DRAM[8478] = 8'b1110011;
DRAM[8479] = 8'b1110011;
DRAM[8480] = 8'b1110010;
DRAM[8481] = 8'b1110010;
DRAM[8482] = 8'b1110010;
DRAM[8483] = 8'b1110011;
DRAM[8484] = 8'b1110011;
DRAM[8485] = 8'b1110100;
DRAM[8486] = 8'b1110100;
DRAM[8487] = 8'b1110100;
DRAM[8488] = 8'b1110101;
DRAM[8489] = 8'b1110110;
DRAM[8490] = 8'b1110110;
DRAM[8491] = 8'b1110111;
DRAM[8492] = 8'b1110111;
DRAM[8493] = 8'b1110110;
DRAM[8494] = 8'b1110110;
DRAM[8495] = 8'b1110101;
DRAM[8496] = 8'b1110101;
DRAM[8497] = 8'b1110110;
DRAM[8498] = 8'b1110111;
DRAM[8499] = 8'b1111000;
DRAM[8500] = 8'b1111000;
DRAM[8501] = 8'b1111000;
DRAM[8502] = 8'b1111000;
DRAM[8503] = 8'b1110111;
DRAM[8504] = 8'b1111000;
DRAM[8505] = 8'b1111001;
DRAM[8506] = 8'b1111001;
DRAM[8507] = 8'b1111010;
DRAM[8508] = 8'b1111010;
DRAM[8509] = 8'b1111001;
DRAM[8510] = 8'b1111001;
DRAM[8511] = 8'b1111000;
DRAM[8512] = 8'b1111010;
DRAM[8513] = 8'b1111010;
DRAM[8514] = 8'b1111010;
DRAM[8515] = 8'b1111010;
DRAM[8516] = 8'b1111010;
DRAM[8517] = 8'b1111010;
DRAM[8518] = 8'b1111010;
DRAM[8519] = 8'b1111010;
DRAM[8520] = 8'b1111101;
DRAM[8521] = 8'b1111101;
DRAM[8522] = 8'b1111100;
DRAM[8523] = 8'b1111100;
DRAM[8524] = 8'b1111011;
DRAM[8525] = 8'b1111011;
DRAM[8526] = 8'b1111011;
DRAM[8527] = 8'b1111011;
DRAM[8528] = 8'b1110111;
DRAM[8529] = 8'b1110111;
DRAM[8530] = 8'b1111000;
DRAM[8531] = 8'b1111010;
DRAM[8532] = 8'b1111100;
DRAM[8533] = 8'b1111101;
DRAM[8534] = 8'b1111101;
DRAM[8535] = 8'b1111100;
DRAM[8536] = 8'b1110111;
DRAM[8537] = 8'b1111111;
DRAM[8538] = 8'b10001001;
DRAM[8539] = 8'b10001000;
DRAM[8540] = 8'b10000011;
DRAM[8541] = 8'b10110101;
DRAM[8542] = 8'b11001101;
DRAM[8543] = 8'b10110011;
DRAM[8544] = 8'b11000100;
DRAM[8545] = 8'b11001101;
DRAM[8546] = 8'b11011101;
DRAM[8547] = 8'b11101101;
DRAM[8548] = 8'b11111001;
DRAM[8549] = 8'b11111111;
DRAM[8550] = 8'b11111111;
DRAM[8551] = 8'b11111111;
DRAM[8552] = 8'b11111011;
DRAM[8553] = 8'b11111011;
DRAM[8554] = 8'b11111011;
DRAM[8555] = 8'b11111011;
DRAM[8556] = 8'b11111011;
DRAM[8557] = 8'b11111011;
DRAM[8558] = 8'b11111011;
DRAM[8559] = 8'b11111011;
DRAM[8560] = 8'b11111001;
DRAM[8561] = 8'b11111010;
DRAM[8562] = 8'b11111010;
DRAM[8563] = 8'b11111011;
DRAM[8564] = 8'b11111100;
DRAM[8565] = 8'b11111101;
DRAM[8566] = 8'b11111110;
DRAM[8567] = 8'b11111110;
DRAM[8568] = 8'b11111110;
DRAM[8569] = 8'b11111110;
DRAM[8570] = 8'b11111110;
DRAM[8571] = 8'b11111111;
DRAM[8572] = 8'b11111111;
DRAM[8573] = 8'b11111111;
DRAM[8574] = 8'b11111111;
DRAM[8575] = 8'b11111111;
DRAM[8576] = 8'b11111111;
DRAM[8577] = 8'b11111111;
DRAM[8578] = 8'b11111111;
DRAM[8579] = 8'b11111111;
DRAM[8580] = 8'b11111111;
DRAM[8581] = 8'b11111111;
DRAM[8582] = 8'b11111111;
DRAM[8583] = 8'b11111111;
DRAM[8584] = 8'b11111111;
DRAM[8585] = 8'b11111111;
DRAM[8586] = 8'b11111111;
DRAM[8587] = 8'b11111111;
DRAM[8588] = 8'b11111111;
DRAM[8589] = 8'b11111111;
DRAM[8590] = 8'b11111111;
DRAM[8591] = 8'b11111111;
DRAM[8592] = 8'b11111111;
DRAM[8593] = 8'b11111111;
DRAM[8594] = 8'b11111111;
DRAM[8595] = 8'b11111111;
DRAM[8596] = 8'b11111111;
DRAM[8597] = 8'b11111111;
DRAM[8598] = 8'b11111111;
DRAM[8599] = 8'b11111111;
DRAM[8600] = 8'b11111100;
DRAM[8601] = 8'b11111100;
DRAM[8602] = 8'b11111101;
DRAM[8603] = 8'b11111101;
DRAM[8604] = 8'b11111101;
DRAM[8605] = 8'b11111110;
DRAM[8606] = 8'b11111110;
DRAM[8607] = 8'b11111110;
DRAM[8608] = 8'b11111100;
DRAM[8609] = 8'b11111100;
DRAM[8610] = 8'b11111100;
DRAM[8611] = 8'b11111100;
DRAM[8612] = 8'b11111100;
DRAM[8613] = 8'b11111100;
DRAM[8614] = 8'b11111100;
DRAM[8615] = 8'b11111100;
DRAM[8616] = 8'b11111111;
DRAM[8617] = 8'b11111100;
DRAM[8618] = 8'b11111000;
DRAM[8619] = 8'b11110101;
DRAM[8620] = 8'b11110100;
DRAM[8621] = 8'b11101100;
DRAM[8622] = 8'b11010101;
DRAM[8623] = 8'b10111110;
DRAM[8624] = 8'b10101001;
DRAM[8625] = 8'b10011111;
DRAM[8626] = 8'b1110100;
DRAM[8627] = 8'b1110010;
DRAM[8628] = 8'b1110000;
DRAM[8629] = 8'b1100110;
DRAM[8630] = 8'b1111001;
DRAM[8631] = 8'b1101111;
DRAM[8632] = 8'b1100101;
DRAM[8633] = 8'b1101100;
DRAM[8634] = 8'b1101110;
DRAM[8635] = 8'b1100111;
DRAM[8636] = 8'b1100000;
DRAM[8637] = 8'b1100100;
DRAM[8638] = 8'b1101111;
DRAM[8639] = 8'b1110111;
DRAM[8640] = 8'b1101110;
DRAM[8641] = 8'b1100001;
DRAM[8642] = 8'b1100100;
DRAM[8643] = 8'b1101110;
DRAM[8644] = 8'b1101110;
DRAM[8645] = 8'b1101101;
DRAM[8646] = 8'b1100110;
DRAM[8647] = 8'b1011000;
DRAM[8648] = 8'b1100101;
DRAM[8649] = 8'b1100011;
DRAM[8650] = 8'b1100000;
DRAM[8651] = 8'b1011111;
DRAM[8652] = 8'b1011111;
DRAM[8653] = 8'b1100000;
DRAM[8654] = 8'b1100000;
DRAM[8655] = 8'b1011111;
DRAM[8656] = 8'b1011101;
DRAM[8657] = 8'b1011101;
DRAM[8658] = 8'b1011100;
DRAM[8659] = 8'b1011100;
DRAM[8660] = 8'b1011011;
DRAM[8661] = 8'b1011010;
DRAM[8662] = 8'b1011001;
DRAM[8663] = 8'b1011001;
DRAM[8664] = 8'b1011001;
DRAM[8665] = 8'b1011001;
DRAM[8666] = 8'b1011000;
DRAM[8667] = 8'b1011000;
DRAM[8668] = 8'b1010111;
DRAM[8669] = 8'b1010110;
DRAM[8670] = 8'b1010101;
DRAM[8671] = 8'b1010101;
DRAM[8672] = 8'b1010100;
DRAM[8673] = 8'b1010100;
DRAM[8674] = 8'b1010100;
DRAM[8675] = 8'b1010100;
DRAM[8676] = 8'b1010100;
DRAM[8677] = 8'b1010100;
DRAM[8678] = 8'b1010100;
DRAM[8679] = 8'b1010100;
DRAM[8680] = 8'b1010001;
DRAM[8681] = 8'b1010010;
DRAM[8682] = 8'b1010010;
DRAM[8683] = 8'b1010011;
DRAM[8684] = 8'b1010011;
DRAM[8685] = 8'b1010010;
DRAM[8686] = 8'b1010010;
DRAM[8687] = 8'b1010001;
DRAM[8688] = 8'b1001111;
DRAM[8689] = 8'b1001111;
DRAM[8690] = 8'b1001111;
DRAM[8691] = 8'b1001110;
DRAM[8692] = 8'b1001110;
DRAM[8693] = 8'b1001110;
DRAM[8694] = 8'b1001101;
DRAM[8695] = 8'b1001101;
DRAM[8696] = 8'b1001101;
DRAM[8697] = 8'b1001101;
DRAM[8698] = 8'b1001101;
DRAM[8699] = 8'b1001100;
DRAM[8700] = 8'b1001100;
DRAM[8701] = 8'b1001100;
DRAM[8702] = 8'b1001011;
DRAM[8703] = 8'b1001011;
DRAM[8704] = 8'b1100001;
DRAM[8705] = 8'b1100010;
DRAM[8706] = 8'b1100100;
DRAM[8707] = 8'b1100101;
DRAM[8708] = 8'b1100110;
DRAM[8709] = 8'b1100111;
DRAM[8710] = 8'b1100111;
DRAM[8711] = 8'b1100111;
DRAM[8712] = 8'b1101000;
DRAM[8713] = 8'b1101000;
DRAM[8714] = 8'b1101000;
DRAM[8715] = 8'b1101001;
DRAM[8716] = 8'b1101001;
DRAM[8717] = 8'b1101010;
DRAM[8718] = 8'b1101010;
DRAM[8719] = 8'b1101010;
DRAM[8720] = 8'b1101011;
DRAM[8721] = 8'b1101011;
DRAM[8722] = 8'b1101100;
DRAM[8723] = 8'b1101101;
DRAM[8724] = 8'b1101101;
DRAM[8725] = 8'b1101110;
DRAM[8726] = 8'b1101111;
DRAM[8727] = 8'b1101111;
DRAM[8728] = 8'b1110001;
DRAM[8729] = 8'b1110001;
DRAM[8730] = 8'b1110001;
DRAM[8731] = 8'b1110001;
DRAM[8732] = 8'b1110010;
DRAM[8733] = 8'b1110010;
DRAM[8734] = 8'b1110010;
DRAM[8735] = 8'b1110011;
DRAM[8736] = 8'b1110010;
DRAM[8737] = 8'b1110010;
DRAM[8738] = 8'b1110010;
DRAM[8739] = 8'b1110011;
DRAM[8740] = 8'b1110011;
DRAM[8741] = 8'b1110100;
DRAM[8742] = 8'b1110100;
DRAM[8743] = 8'b1110100;
DRAM[8744] = 8'b1110101;
DRAM[8745] = 8'b1110101;
DRAM[8746] = 8'b1110110;
DRAM[8747] = 8'b1110111;
DRAM[8748] = 8'b1110111;
DRAM[8749] = 8'b1110110;
DRAM[8750] = 8'b1110110;
DRAM[8751] = 8'b1110101;
DRAM[8752] = 8'b1110110;
DRAM[8753] = 8'b1110111;
DRAM[8754] = 8'b1111000;
DRAM[8755] = 8'b1111000;
DRAM[8756] = 8'b1111001;
DRAM[8757] = 8'b1111001;
DRAM[8758] = 8'b1111000;
DRAM[8759] = 8'b1111000;
DRAM[8760] = 8'b1111001;
DRAM[8761] = 8'b1111001;
DRAM[8762] = 8'b1111010;
DRAM[8763] = 8'b1111010;
DRAM[8764] = 8'b1111010;
DRAM[8765] = 8'b1111010;
DRAM[8766] = 8'b1111001;
DRAM[8767] = 8'b1111001;
DRAM[8768] = 8'b1111010;
DRAM[8769] = 8'b1111010;
DRAM[8770] = 8'b1111010;
DRAM[8771] = 8'b1111010;
DRAM[8772] = 8'b1111010;
DRAM[8773] = 8'b1111010;
DRAM[8774] = 8'b1111010;
DRAM[8775] = 8'b1111010;
DRAM[8776] = 8'b1111101;
DRAM[8777] = 8'b1111100;
DRAM[8778] = 8'b1111100;
DRAM[8779] = 8'b1111100;
DRAM[8780] = 8'b1111100;
DRAM[8781] = 8'b1111011;
DRAM[8782] = 8'b1111011;
DRAM[8783] = 8'b1111011;
DRAM[8784] = 8'b1110111;
DRAM[8785] = 8'b1111000;
DRAM[8786] = 8'b1111010;
DRAM[8787] = 8'b1111011;
DRAM[8788] = 8'b1111100;
DRAM[8789] = 8'b1111101;
DRAM[8790] = 8'b1111101;
DRAM[8791] = 8'b1111101;
DRAM[8792] = 8'b10001100;
DRAM[8793] = 8'b1110011;
DRAM[8794] = 8'b10000001;
DRAM[8795] = 8'b10001000;
DRAM[8796] = 8'b10000111;
DRAM[8797] = 8'b10100000;
DRAM[8798] = 8'b11011101;
DRAM[8799] = 8'b11110111;
DRAM[8800] = 8'b11101110;
DRAM[8801] = 8'b11110100;
DRAM[8802] = 8'b11111101;
DRAM[8803] = 8'b11111111;
DRAM[8804] = 8'b11111111;
DRAM[8805] = 8'b11111111;
DRAM[8806] = 8'b11111010;
DRAM[8807] = 8'b11110101;
DRAM[8808] = 8'b11111110;
DRAM[8809] = 8'b11111110;
DRAM[8810] = 8'b11111110;
DRAM[8811] = 8'b11111110;
DRAM[8812] = 8'b11111110;
DRAM[8813] = 8'b11111110;
DRAM[8814] = 8'b11111110;
DRAM[8815] = 8'b11111110;
DRAM[8816] = 8'b11111011;
DRAM[8817] = 8'b11111011;
DRAM[8818] = 8'b11111100;
DRAM[8819] = 8'b11111101;
DRAM[8820] = 8'b11111101;
DRAM[8821] = 8'b11111110;
DRAM[8822] = 8'b11111110;
DRAM[8823] = 8'b11111111;
DRAM[8824] = 8'b11111110;
DRAM[8825] = 8'b11111110;
DRAM[8826] = 8'b11111110;
DRAM[8827] = 8'b11111111;
DRAM[8828] = 8'b11111111;
DRAM[8829] = 8'b11111111;
DRAM[8830] = 8'b11111111;
DRAM[8831] = 8'b11111111;
DRAM[8832] = 8'b11111111;
DRAM[8833] = 8'b11111111;
DRAM[8834] = 8'b11111111;
DRAM[8835] = 8'b11111111;
DRAM[8836] = 8'b11111111;
DRAM[8837] = 8'b11111111;
DRAM[8838] = 8'b11111111;
DRAM[8839] = 8'b11111111;
DRAM[8840] = 8'b11111111;
DRAM[8841] = 8'b11111111;
DRAM[8842] = 8'b11111111;
DRAM[8843] = 8'b11111111;
DRAM[8844] = 8'b11111111;
DRAM[8845] = 8'b11111111;
DRAM[8846] = 8'b11111111;
DRAM[8847] = 8'b11111111;
DRAM[8848] = 8'b11111111;
DRAM[8849] = 8'b11111111;
DRAM[8850] = 8'b11111111;
DRAM[8851] = 8'b11111111;
DRAM[8852] = 8'b11111111;
DRAM[8853] = 8'b11111111;
DRAM[8854] = 8'b11111111;
DRAM[8855] = 8'b11111111;
DRAM[8856] = 8'b11111100;
DRAM[8857] = 8'b11111101;
DRAM[8858] = 8'b11111101;
DRAM[8859] = 8'b11111101;
DRAM[8860] = 8'b11111110;
DRAM[8861] = 8'b11111110;
DRAM[8862] = 8'b11111110;
DRAM[8863] = 8'b11111110;
DRAM[8864] = 8'b11111110;
DRAM[8865] = 8'b11111110;
DRAM[8866] = 8'b11111110;
DRAM[8867] = 8'b11111110;
DRAM[8868] = 8'b11111110;
DRAM[8869] = 8'b11111110;
DRAM[8870] = 8'b11111110;
DRAM[8871] = 8'b11111110;
DRAM[8872] = 8'b11111000;
DRAM[8873] = 8'b11111101;
DRAM[8874] = 8'b11111111;
DRAM[8875] = 8'b11111111;
DRAM[8876] = 8'b11111101;
DRAM[8877] = 8'b11111001;
DRAM[8878] = 8'b11110010;
DRAM[8879] = 8'b11101011;
DRAM[8880] = 8'b11011000;
DRAM[8881] = 8'b10101010;
DRAM[8882] = 8'b1101010;
DRAM[8883] = 8'b1111000;
DRAM[8884] = 8'b10000111;
DRAM[8885] = 8'b1110110;
DRAM[8886] = 8'b1111010;
DRAM[8887] = 8'b1101010;
DRAM[8888] = 8'b1110010;
DRAM[8889] = 8'b1111000;
DRAM[8890] = 8'b1110110;
DRAM[8891] = 8'b1101110;
DRAM[8892] = 8'b1110000;
DRAM[8893] = 8'b1111001;
DRAM[8894] = 8'b1111001;
DRAM[8895] = 8'b1101111;
DRAM[8896] = 8'b1101010;
DRAM[8897] = 8'b1100010;
DRAM[8898] = 8'b1100101;
DRAM[8899] = 8'b1101010;
DRAM[8900] = 8'b1100101;
DRAM[8901] = 8'b1100101;
DRAM[8902] = 8'b1100110;
DRAM[8903] = 8'b1011111;
DRAM[8904] = 8'b1100110;
DRAM[8905] = 8'b1100100;
DRAM[8906] = 8'b1100001;
DRAM[8907] = 8'b1100001;
DRAM[8908] = 8'b1100010;
DRAM[8909] = 8'b1100010;
DRAM[8910] = 8'b1100001;
DRAM[8911] = 8'b1100000;
DRAM[8912] = 8'b1011101;
DRAM[8913] = 8'b1011101;
DRAM[8914] = 8'b1011101;
DRAM[8915] = 8'b1011100;
DRAM[8916] = 8'b1011011;
DRAM[8917] = 8'b1011010;
DRAM[8918] = 8'b1011010;
DRAM[8919] = 8'b1011001;
DRAM[8920] = 8'b1011001;
DRAM[8921] = 8'b1011001;
DRAM[8922] = 8'b1011001;
DRAM[8923] = 8'b1011000;
DRAM[8924] = 8'b1010111;
DRAM[8925] = 8'b1010110;
DRAM[8926] = 8'b1010110;
DRAM[8927] = 8'b1010101;
DRAM[8928] = 8'b1010100;
DRAM[8929] = 8'b1010100;
DRAM[8930] = 8'b1010100;
DRAM[8931] = 8'b1010100;
DRAM[8932] = 8'b1010100;
DRAM[8933] = 8'b1010100;
DRAM[8934] = 8'b1010100;
DRAM[8935] = 8'b1010100;
DRAM[8936] = 8'b1010001;
DRAM[8937] = 8'b1010010;
DRAM[8938] = 8'b1010010;
DRAM[8939] = 8'b1010011;
DRAM[8940] = 8'b1010011;
DRAM[8941] = 8'b1010010;
DRAM[8942] = 8'b1010010;
DRAM[8943] = 8'b1010001;
DRAM[8944] = 8'b1001111;
DRAM[8945] = 8'b1001111;
DRAM[8946] = 8'b1001111;
DRAM[8947] = 8'b1001111;
DRAM[8948] = 8'b1001110;
DRAM[8949] = 8'b1001110;
DRAM[8950] = 8'b1001110;
DRAM[8951] = 8'b1001101;
DRAM[8952] = 8'b1001101;
DRAM[8953] = 8'b1001101;
DRAM[8954] = 8'b1001101;
DRAM[8955] = 8'b1001101;
DRAM[8956] = 8'b1001100;
DRAM[8957] = 8'b1001100;
DRAM[8958] = 8'b1001100;
DRAM[8959] = 8'b1001011;
DRAM[8960] = 8'b1100010;
DRAM[8961] = 8'b1100011;
DRAM[8962] = 8'b1100100;
DRAM[8963] = 8'b1100101;
DRAM[8964] = 8'b1100110;
DRAM[8965] = 8'b1100111;
DRAM[8966] = 8'b1100111;
DRAM[8967] = 8'b1100111;
DRAM[8968] = 8'b1101000;
DRAM[8969] = 8'b1101000;
DRAM[8970] = 8'b1101000;
DRAM[8971] = 8'b1101001;
DRAM[8972] = 8'b1101001;
DRAM[8973] = 8'b1101010;
DRAM[8974] = 8'b1101010;
DRAM[8975] = 8'b1101010;
DRAM[8976] = 8'b1101011;
DRAM[8977] = 8'b1101011;
DRAM[8978] = 8'b1101100;
DRAM[8979] = 8'b1101101;
DRAM[8980] = 8'b1101101;
DRAM[8981] = 8'b1101110;
DRAM[8982] = 8'b1101111;
DRAM[8983] = 8'b1101111;
DRAM[8984] = 8'b1110000;
DRAM[8985] = 8'b1110000;
DRAM[8986] = 8'b1110001;
DRAM[8987] = 8'b1110001;
DRAM[8988] = 8'b1110001;
DRAM[8989] = 8'b1110010;
DRAM[8990] = 8'b1110010;
DRAM[8991] = 8'b1110010;
DRAM[8992] = 8'b1110010;
DRAM[8993] = 8'b1110010;
DRAM[8994] = 8'b1110010;
DRAM[8995] = 8'b1110011;
DRAM[8996] = 8'b1110011;
DRAM[8997] = 8'b1110100;
DRAM[8998] = 8'b1110100;
DRAM[8999] = 8'b1110100;
DRAM[9000] = 8'b1110100;
DRAM[9001] = 8'b1110101;
DRAM[9002] = 8'b1110110;
DRAM[9003] = 8'b1110111;
DRAM[9004] = 8'b1110111;
DRAM[9005] = 8'b1110111;
DRAM[9006] = 8'b1110110;
DRAM[9007] = 8'b1110110;
DRAM[9008] = 8'b1110111;
DRAM[9009] = 8'b1110111;
DRAM[9010] = 8'b1111000;
DRAM[9011] = 8'b1111001;
DRAM[9012] = 8'b1111010;
DRAM[9013] = 8'b1111010;
DRAM[9014] = 8'b1111001;
DRAM[9015] = 8'b1111001;
DRAM[9016] = 8'b1111001;
DRAM[9017] = 8'b1111001;
DRAM[9018] = 8'b1111010;
DRAM[9019] = 8'b1111011;
DRAM[9020] = 8'b1111011;
DRAM[9021] = 8'b1111010;
DRAM[9022] = 8'b1111001;
DRAM[9023] = 8'b1111001;
DRAM[9024] = 8'b1111011;
DRAM[9025] = 8'b1111011;
DRAM[9026] = 8'b1111011;
DRAM[9027] = 8'b1111011;
DRAM[9028] = 8'b1111011;
DRAM[9029] = 8'b1111011;
DRAM[9030] = 8'b1111011;
DRAM[9031] = 8'b1111011;
DRAM[9032] = 8'b1111011;
DRAM[9033] = 8'b1111011;
DRAM[9034] = 8'b1111011;
DRAM[9035] = 8'b1111011;
DRAM[9036] = 8'b1111010;
DRAM[9037] = 8'b1111010;
DRAM[9038] = 8'b1111010;
DRAM[9039] = 8'b1111010;
DRAM[9040] = 8'b1111011;
DRAM[9041] = 8'b1111101;
DRAM[9042] = 8'b1111110;
DRAM[9043] = 8'b1111110;
DRAM[9044] = 8'b1111101;
DRAM[9045] = 8'b1111100;
DRAM[9046] = 8'b1111100;
DRAM[9047] = 8'b1111101;
DRAM[9048] = 8'b1111001;
DRAM[9049] = 8'b10100110;
DRAM[9050] = 8'b10101101;
DRAM[9051] = 8'b10000111;
DRAM[9052] = 8'b10101101;
DRAM[9053] = 8'b11001100;
DRAM[9054] = 8'b11101111;
DRAM[9055] = 8'b11111100;
DRAM[9056] = 8'b11111101;
DRAM[9057] = 8'b11111101;
DRAM[9058] = 8'b11111101;
DRAM[9059] = 8'b11111101;
DRAM[9060] = 8'b11111100;
DRAM[9061] = 8'b11111100;
DRAM[9062] = 8'b11111011;
DRAM[9063] = 8'b11111010;
DRAM[9064] = 8'b11111110;
DRAM[9065] = 8'b11111110;
DRAM[9066] = 8'b11111110;
DRAM[9067] = 8'b11111110;
DRAM[9068] = 8'b11111110;
DRAM[9069] = 8'b11111110;
DRAM[9070] = 8'b11111110;
DRAM[9071] = 8'b11111110;
DRAM[9072] = 8'b11111101;
DRAM[9073] = 8'b11111101;
DRAM[9074] = 8'b11111101;
DRAM[9075] = 8'b11111110;
DRAM[9076] = 8'b11111110;
DRAM[9077] = 8'b11111111;
DRAM[9078] = 8'b11111111;
DRAM[9079] = 8'b11111111;
DRAM[9080] = 8'b11111110;
DRAM[9081] = 8'b11111110;
DRAM[9082] = 8'b11111110;
DRAM[9083] = 8'b11111111;
DRAM[9084] = 8'b11111111;
DRAM[9085] = 8'b11111111;
DRAM[9086] = 8'b11111111;
DRAM[9087] = 8'b11111111;
DRAM[9088] = 8'b11111111;
DRAM[9089] = 8'b11111111;
DRAM[9090] = 8'b11111111;
DRAM[9091] = 8'b11111111;
DRAM[9092] = 8'b11111111;
DRAM[9093] = 8'b11111111;
DRAM[9094] = 8'b11111111;
DRAM[9095] = 8'b11111111;
DRAM[9096] = 8'b11111111;
DRAM[9097] = 8'b11111111;
DRAM[9098] = 8'b11111111;
DRAM[9099] = 8'b11111111;
DRAM[9100] = 8'b11111111;
DRAM[9101] = 8'b11111111;
DRAM[9102] = 8'b11111111;
DRAM[9103] = 8'b11111111;
DRAM[9104] = 8'b11111111;
DRAM[9105] = 8'b11111111;
DRAM[9106] = 8'b11111111;
DRAM[9107] = 8'b11111111;
DRAM[9108] = 8'b11111111;
DRAM[9109] = 8'b11111111;
DRAM[9110] = 8'b11111111;
DRAM[9111] = 8'b11111111;
DRAM[9112] = 8'b11111101;
DRAM[9113] = 8'b11111101;
DRAM[9114] = 8'b11111101;
DRAM[9115] = 8'b11111110;
DRAM[9116] = 8'b11111110;
DRAM[9117] = 8'b11111110;
DRAM[9118] = 8'b11111111;
DRAM[9119] = 8'b11111111;
DRAM[9120] = 8'b11111111;
DRAM[9121] = 8'b11111111;
DRAM[9122] = 8'b11111111;
DRAM[9123] = 8'b11111111;
DRAM[9124] = 8'b11111111;
DRAM[9125] = 8'b11111111;
DRAM[9126] = 8'b11111111;
DRAM[9127] = 8'b11111111;
DRAM[9128] = 8'b11110110;
DRAM[9129] = 8'b11111100;
DRAM[9130] = 8'b11111111;
DRAM[9131] = 8'b11111111;
DRAM[9132] = 8'b11111010;
DRAM[9133] = 8'b11111000;
DRAM[9134] = 8'b11111001;
DRAM[9135] = 8'b11111011;
DRAM[9136] = 8'b11110001;
DRAM[9137] = 8'b10110101;
DRAM[9138] = 8'b10011101;
DRAM[9139] = 8'b10001011;
DRAM[9140] = 8'b10001011;
DRAM[9141] = 8'b10001010;
DRAM[9142] = 8'b1101111;
DRAM[9143] = 8'b1111101;
DRAM[9144] = 8'b10011001;
DRAM[9145] = 8'b10000000;
DRAM[9146] = 8'b1101000;
DRAM[9147] = 8'b1101011;
DRAM[9148] = 8'b10000110;
DRAM[9149] = 8'b10011011;
DRAM[9150] = 8'b10010010;
DRAM[9151] = 8'b1111110;
DRAM[9152] = 8'b1100000;
DRAM[9153] = 8'b1101101;
DRAM[9154] = 8'b1111010;
DRAM[9155] = 8'b1110000;
DRAM[9156] = 8'b1011011;
DRAM[9157] = 8'b1011110;
DRAM[9158] = 8'b1101001;
DRAM[9159] = 8'b1100111;
DRAM[9160] = 8'b1100110;
DRAM[9161] = 8'b1100100;
DRAM[9162] = 8'b1100010;
DRAM[9163] = 8'b1100010;
DRAM[9164] = 8'b1100010;
DRAM[9165] = 8'b1100010;
DRAM[9166] = 8'b1100001;
DRAM[9167] = 8'b1011111;
DRAM[9168] = 8'b1011110;
DRAM[9169] = 8'b1011110;
DRAM[9170] = 8'b1011101;
DRAM[9171] = 8'b1011100;
DRAM[9172] = 8'b1011011;
DRAM[9173] = 8'b1011011;
DRAM[9174] = 8'b1011010;
DRAM[9175] = 8'b1011010;
DRAM[9176] = 8'b1011010;
DRAM[9177] = 8'b1011010;
DRAM[9178] = 8'b1011001;
DRAM[9179] = 8'b1011000;
DRAM[9180] = 8'b1010111;
DRAM[9181] = 8'b1010111;
DRAM[9182] = 8'b1010110;
DRAM[9183] = 8'b1010110;
DRAM[9184] = 8'b1010100;
DRAM[9185] = 8'b1010100;
DRAM[9186] = 8'b1010100;
DRAM[9187] = 8'b1010100;
DRAM[9188] = 8'b1010100;
DRAM[9189] = 8'b1010100;
DRAM[9190] = 8'b1010100;
DRAM[9191] = 8'b1010100;
DRAM[9192] = 8'b1010001;
DRAM[9193] = 8'b1010010;
DRAM[9194] = 8'b1010010;
DRAM[9195] = 8'b1010011;
DRAM[9196] = 8'b1010011;
DRAM[9197] = 8'b1010010;
DRAM[9198] = 8'b1010010;
DRAM[9199] = 8'b1010001;
DRAM[9200] = 8'b1010000;
DRAM[9201] = 8'b1010000;
DRAM[9202] = 8'b1001111;
DRAM[9203] = 8'b1001111;
DRAM[9204] = 8'b1001111;
DRAM[9205] = 8'b1001110;
DRAM[9206] = 8'b1001110;
DRAM[9207] = 8'b1001110;
DRAM[9208] = 8'b1001110;
DRAM[9209] = 8'b1001110;
DRAM[9210] = 8'b1001101;
DRAM[9211] = 8'b1001101;
DRAM[9212] = 8'b1001101;
DRAM[9213] = 8'b1001100;
DRAM[9214] = 8'b1001100;
DRAM[9215] = 8'b1001100;
DRAM[9216] = 8'b1100010;
DRAM[9217] = 8'b1100011;
DRAM[9218] = 8'b1100100;
DRAM[9219] = 8'b1100101;
DRAM[9220] = 8'b1100110;
DRAM[9221] = 8'b1100110;
DRAM[9222] = 8'b1100110;
DRAM[9223] = 8'b1100110;
DRAM[9224] = 8'b1101000;
DRAM[9225] = 8'b1101000;
DRAM[9226] = 8'b1101000;
DRAM[9227] = 8'b1101001;
DRAM[9228] = 8'b1101001;
DRAM[9229] = 8'b1101010;
DRAM[9230] = 8'b1101010;
DRAM[9231] = 8'b1101010;
DRAM[9232] = 8'b1101011;
DRAM[9233] = 8'b1101011;
DRAM[9234] = 8'b1101100;
DRAM[9235] = 8'b1101101;
DRAM[9236] = 8'b1101101;
DRAM[9237] = 8'b1101110;
DRAM[9238] = 8'b1101111;
DRAM[9239] = 8'b1101111;
DRAM[9240] = 8'b1110000;
DRAM[9241] = 8'b1110000;
DRAM[9242] = 8'b1110000;
DRAM[9243] = 8'b1110001;
DRAM[9244] = 8'b1110001;
DRAM[9245] = 8'b1110001;
DRAM[9246] = 8'b1110010;
DRAM[9247] = 8'b1110010;
DRAM[9248] = 8'b1110010;
DRAM[9249] = 8'b1110010;
DRAM[9250] = 8'b1110010;
DRAM[9251] = 8'b1110011;
DRAM[9252] = 8'b1110011;
DRAM[9253] = 8'b1110100;
DRAM[9254] = 8'b1110100;
DRAM[9255] = 8'b1110100;
DRAM[9256] = 8'b1110100;
DRAM[9257] = 8'b1110101;
DRAM[9258] = 8'b1110110;
DRAM[9259] = 8'b1110111;
DRAM[9260] = 8'b1110111;
DRAM[9261] = 8'b1110111;
DRAM[9262] = 8'b1110111;
DRAM[9263] = 8'b1110111;
DRAM[9264] = 8'b1111000;
DRAM[9265] = 8'b1111000;
DRAM[9266] = 8'b1111001;
DRAM[9267] = 8'b1111010;
DRAM[9268] = 8'b1111010;
DRAM[9269] = 8'b1111010;
DRAM[9270] = 8'b1111010;
DRAM[9271] = 8'b1111010;
DRAM[9272] = 8'b1111001;
DRAM[9273] = 8'b1111010;
DRAM[9274] = 8'b1111011;
DRAM[9275] = 8'b1111011;
DRAM[9276] = 8'b1111011;
DRAM[9277] = 8'b1111011;
DRAM[9278] = 8'b1111010;
DRAM[9279] = 8'b1111001;
DRAM[9280] = 8'b1111011;
DRAM[9281] = 8'b1111011;
DRAM[9282] = 8'b1111011;
DRAM[9283] = 8'b1111011;
DRAM[9284] = 8'b1111011;
DRAM[9285] = 8'b1111011;
DRAM[9286] = 8'b1111011;
DRAM[9287] = 8'b1111011;
DRAM[9288] = 8'b1111001;
DRAM[9289] = 8'b1111001;
DRAM[9290] = 8'b1111001;
DRAM[9291] = 8'b1111001;
DRAM[9292] = 8'b1111001;
DRAM[9293] = 8'b1111001;
DRAM[9294] = 8'b1111001;
DRAM[9295] = 8'b1111001;
DRAM[9296] = 8'b1111101;
DRAM[9297] = 8'b1111110;
DRAM[9298] = 8'b10000000;
DRAM[9299] = 8'b1111111;
DRAM[9300] = 8'b1111110;
DRAM[9301] = 8'b1111110;
DRAM[9302] = 8'b10000000;
DRAM[9303] = 8'b10000011;
DRAM[9304] = 8'b1110001;
DRAM[9305] = 8'b10011110;
DRAM[9306] = 8'b10111111;
DRAM[9307] = 8'b11000010;
DRAM[9308] = 8'b11110011;
DRAM[9309] = 8'b11110111;
DRAM[9310] = 8'b11111000;
DRAM[9311] = 8'b11111000;
DRAM[9312] = 8'b11111111;
DRAM[9313] = 8'b11111101;
DRAM[9314] = 8'b11111011;
DRAM[9315] = 8'b11111010;
DRAM[9316] = 8'b11111011;
DRAM[9317] = 8'b11111110;
DRAM[9318] = 8'b11111111;
DRAM[9319] = 8'b11111111;
DRAM[9320] = 8'b11111110;
DRAM[9321] = 8'b11111110;
DRAM[9322] = 8'b11111110;
DRAM[9323] = 8'b11111110;
DRAM[9324] = 8'b11111110;
DRAM[9325] = 8'b11111110;
DRAM[9326] = 8'b11111110;
DRAM[9327] = 8'b11111110;
DRAM[9328] = 8'b11111110;
DRAM[9329] = 8'b11111110;
DRAM[9330] = 8'b11111110;
DRAM[9331] = 8'b11111110;
DRAM[9332] = 8'b11111110;
DRAM[9333] = 8'b11111111;
DRAM[9334] = 8'b11111111;
DRAM[9335] = 8'b11111111;
DRAM[9336] = 8'b11111110;
DRAM[9337] = 8'b11111110;
DRAM[9338] = 8'b11111110;
DRAM[9339] = 8'b11111111;
DRAM[9340] = 8'b11111111;
DRAM[9341] = 8'b11111111;
DRAM[9342] = 8'b11111111;
DRAM[9343] = 8'b11111111;
DRAM[9344] = 8'b11111111;
DRAM[9345] = 8'b11111111;
DRAM[9346] = 8'b11111111;
DRAM[9347] = 8'b11111111;
DRAM[9348] = 8'b11111111;
DRAM[9349] = 8'b11111111;
DRAM[9350] = 8'b11111111;
DRAM[9351] = 8'b11111111;
DRAM[9352] = 8'b11111111;
DRAM[9353] = 8'b11111111;
DRAM[9354] = 8'b11111111;
DRAM[9355] = 8'b11111111;
DRAM[9356] = 8'b11111111;
DRAM[9357] = 8'b11111111;
DRAM[9358] = 8'b11111111;
DRAM[9359] = 8'b11111111;
DRAM[9360] = 8'b11111111;
DRAM[9361] = 8'b11111111;
DRAM[9362] = 8'b11111111;
DRAM[9363] = 8'b11111111;
DRAM[9364] = 8'b11111111;
DRAM[9365] = 8'b11111111;
DRAM[9366] = 8'b11111111;
DRAM[9367] = 8'b11111111;
DRAM[9368] = 8'b11111101;
DRAM[9369] = 8'b11111101;
DRAM[9370] = 8'b11111110;
DRAM[9371] = 8'b11111110;
DRAM[9372] = 8'b11111110;
DRAM[9373] = 8'b11111111;
DRAM[9374] = 8'b11111111;
DRAM[9375] = 8'b11111111;
DRAM[9376] = 8'b11111110;
DRAM[9377] = 8'b11111110;
DRAM[9378] = 8'b11111110;
DRAM[9379] = 8'b11111110;
DRAM[9380] = 8'b11111110;
DRAM[9381] = 8'b11111110;
DRAM[9382] = 8'b11111110;
DRAM[9383] = 8'b11111110;
DRAM[9384] = 8'b11111110;
DRAM[9385] = 8'b11111111;
DRAM[9386] = 8'b11111111;
DRAM[9387] = 8'b11111110;
DRAM[9388] = 8'b11111100;
DRAM[9389] = 8'b11111010;
DRAM[9390] = 8'b11111011;
DRAM[9391] = 8'b11111110;
DRAM[9392] = 8'b11111011;
DRAM[9393] = 8'b11100010;
DRAM[9394] = 8'b11011100;
DRAM[9395] = 8'b10110001;
DRAM[9396] = 8'b10010000;
DRAM[9397] = 8'b10001101;
DRAM[9398] = 8'b10001001;
DRAM[9399] = 8'b10101010;
DRAM[9400] = 8'b10001001;
DRAM[9401] = 8'b1111110;
DRAM[9402] = 8'b10000110;
DRAM[9403] = 8'b10100101;
DRAM[9404] = 8'b10111011;
DRAM[9405] = 8'b10101110;
DRAM[9406] = 8'b10010000;
DRAM[9407] = 8'b1111011;
DRAM[9408] = 8'b1101111;
DRAM[9409] = 8'b10000010;
DRAM[9410] = 8'b10001110;
DRAM[9411] = 8'b1111101;
DRAM[9412] = 8'b1100111;
DRAM[9413] = 8'b1101010;
DRAM[9414] = 8'b1101101;
DRAM[9415] = 8'b1011111;
DRAM[9416] = 8'b1100101;
DRAM[9417] = 8'b1100011;
DRAM[9418] = 8'b1100010;
DRAM[9419] = 8'b1100010;
DRAM[9420] = 8'b1100010;
DRAM[9421] = 8'b1100010;
DRAM[9422] = 8'b1100000;
DRAM[9423] = 8'b1011110;
DRAM[9424] = 8'b1011110;
DRAM[9425] = 8'b1011110;
DRAM[9426] = 8'b1011101;
DRAM[9427] = 8'b1011101;
DRAM[9428] = 8'b1011100;
DRAM[9429] = 8'b1011011;
DRAM[9430] = 8'b1011010;
DRAM[9431] = 8'b1011010;
DRAM[9432] = 8'b1011010;
DRAM[9433] = 8'b1011010;
DRAM[9434] = 8'b1011001;
DRAM[9435] = 8'b1011001;
DRAM[9436] = 8'b1011000;
DRAM[9437] = 8'b1010111;
DRAM[9438] = 8'b1010110;
DRAM[9439] = 8'b1010110;
DRAM[9440] = 8'b1010100;
DRAM[9441] = 8'b1010100;
DRAM[9442] = 8'b1010100;
DRAM[9443] = 8'b1010100;
DRAM[9444] = 8'b1010100;
DRAM[9445] = 8'b1010100;
DRAM[9446] = 8'b1010100;
DRAM[9447] = 8'b1010100;
DRAM[9448] = 8'b1010001;
DRAM[9449] = 8'b1010010;
DRAM[9450] = 8'b1010010;
DRAM[9451] = 8'b1010011;
DRAM[9452] = 8'b1010011;
DRAM[9453] = 8'b1010010;
DRAM[9454] = 8'b1010010;
DRAM[9455] = 8'b1010001;
DRAM[9456] = 8'b1010000;
DRAM[9457] = 8'b1010000;
DRAM[9458] = 8'b1010000;
DRAM[9459] = 8'b1001111;
DRAM[9460] = 8'b1001111;
DRAM[9461] = 8'b1001111;
DRAM[9462] = 8'b1001110;
DRAM[9463] = 8'b1001110;
DRAM[9464] = 8'b1001110;
DRAM[9465] = 8'b1001110;
DRAM[9466] = 8'b1001110;
DRAM[9467] = 8'b1001101;
DRAM[9468] = 8'b1001101;
DRAM[9469] = 8'b1001101;
DRAM[9470] = 8'b1001100;
DRAM[9471] = 8'b1001100;
DRAM[9472] = 8'b1100011;
DRAM[9473] = 8'b1100100;
DRAM[9474] = 8'b1100101;
DRAM[9475] = 8'b1100110;
DRAM[9476] = 8'b1100110;
DRAM[9477] = 8'b1100110;
DRAM[9478] = 8'b1100110;
DRAM[9479] = 8'b1100101;
DRAM[9480] = 8'b1101000;
DRAM[9481] = 8'b1101000;
DRAM[9482] = 8'b1101000;
DRAM[9483] = 8'b1101001;
DRAM[9484] = 8'b1101001;
DRAM[9485] = 8'b1101010;
DRAM[9486] = 8'b1101010;
DRAM[9487] = 8'b1101010;
DRAM[9488] = 8'b1101011;
DRAM[9489] = 8'b1101011;
DRAM[9490] = 8'b1101100;
DRAM[9491] = 8'b1101101;
DRAM[9492] = 8'b1101101;
DRAM[9493] = 8'b1101110;
DRAM[9494] = 8'b1101111;
DRAM[9495] = 8'b1101111;
DRAM[9496] = 8'b1101111;
DRAM[9497] = 8'b1110000;
DRAM[9498] = 8'b1110000;
DRAM[9499] = 8'b1110000;
DRAM[9500] = 8'b1110001;
DRAM[9501] = 8'b1110001;
DRAM[9502] = 8'b1110001;
DRAM[9503] = 8'b1110001;
DRAM[9504] = 8'b1110010;
DRAM[9505] = 8'b1110010;
DRAM[9506] = 8'b1110010;
DRAM[9507] = 8'b1110011;
DRAM[9508] = 8'b1110011;
DRAM[9509] = 8'b1110100;
DRAM[9510] = 8'b1110100;
DRAM[9511] = 8'b1110100;
DRAM[9512] = 8'b1110011;
DRAM[9513] = 8'b1110100;
DRAM[9514] = 8'b1110101;
DRAM[9515] = 8'b1110110;
DRAM[9516] = 8'b1110111;
DRAM[9517] = 8'b1110111;
DRAM[9518] = 8'b1110111;
DRAM[9519] = 8'b1110111;
DRAM[9520] = 8'b1111000;
DRAM[9521] = 8'b1111001;
DRAM[9522] = 8'b1111010;
DRAM[9523] = 8'b1111011;
DRAM[9524] = 8'b1111011;
DRAM[9525] = 8'b1111011;
DRAM[9526] = 8'b1111011;
DRAM[9527] = 8'b1111010;
DRAM[9528] = 8'b1111010;
DRAM[9529] = 8'b1111010;
DRAM[9530] = 8'b1111011;
DRAM[9531] = 8'b1111011;
DRAM[9532] = 8'b1111011;
DRAM[9533] = 8'b1111011;
DRAM[9534] = 8'b1111010;
DRAM[9535] = 8'b1111010;
DRAM[9536] = 8'b1111100;
DRAM[9537] = 8'b1111100;
DRAM[9538] = 8'b1111100;
DRAM[9539] = 8'b1111100;
DRAM[9540] = 8'b1111100;
DRAM[9541] = 8'b1111100;
DRAM[9542] = 8'b1111100;
DRAM[9543] = 8'b1111100;
DRAM[9544] = 8'b1111000;
DRAM[9545] = 8'b1111001;
DRAM[9546] = 8'b1111001;
DRAM[9547] = 8'b1111001;
DRAM[9548] = 8'b1111001;
DRAM[9549] = 8'b1111010;
DRAM[9550] = 8'b1111010;
DRAM[9551] = 8'b1111010;
DRAM[9552] = 8'b1111011;
DRAM[9553] = 8'b1111101;
DRAM[9554] = 8'b1111111;
DRAM[9555] = 8'b1111111;
DRAM[9556] = 8'b1111111;
DRAM[9557] = 8'b10000011;
DRAM[9558] = 8'b10001001;
DRAM[9559] = 8'b10001111;
DRAM[9560] = 8'b10011111;
DRAM[9561] = 8'b1111101;
DRAM[9562] = 8'b10101101;
DRAM[9563] = 8'b11110111;
DRAM[9564] = 8'b11111111;
DRAM[9565] = 8'b11101010;
DRAM[9566] = 8'b11110100;
DRAM[9567] = 8'b11111111;
DRAM[9568] = 8'b11111011;
DRAM[9569] = 8'b11111011;
DRAM[9570] = 8'b11111100;
DRAM[9571] = 8'b11111100;
DRAM[9572] = 8'b11111100;
DRAM[9573] = 8'b11111100;
DRAM[9574] = 8'b11111100;
DRAM[9575] = 8'b11111100;
DRAM[9576] = 8'b11111101;
DRAM[9577] = 8'b11111101;
DRAM[9578] = 8'b11111101;
DRAM[9579] = 8'b11111101;
DRAM[9580] = 8'b11111101;
DRAM[9581] = 8'b11111101;
DRAM[9582] = 8'b11111101;
DRAM[9583] = 8'b11111101;
DRAM[9584] = 8'b11111110;
DRAM[9585] = 8'b11111110;
DRAM[9586] = 8'b11111110;
DRAM[9587] = 8'b11111110;
DRAM[9588] = 8'b11111110;
DRAM[9589] = 8'b11111110;
DRAM[9590] = 8'b11111110;
DRAM[9591] = 8'b11111110;
DRAM[9592] = 8'b11111110;
DRAM[9593] = 8'b11111110;
DRAM[9594] = 8'b11111110;
DRAM[9595] = 8'b11111111;
DRAM[9596] = 8'b11111111;
DRAM[9597] = 8'b11111111;
DRAM[9598] = 8'b11111111;
DRAM[9599] = 8'b11111111;
DRAM[9600] = 8'b11111111;
DRAM[9601] = 8'b11111111;
DRAM[9602] = 8'b11111111;
DRAM[9603] = 8'b11111111;
DRAM[9604] = 8'b11111111;
DRAM[9605] = 8'b11111111;
DRAM[9606] = 8'b11111111;
DRAM[9607] = 8'b11111111;
DRAM[9608] = 8'b11111111;
DRAM[9609] = 8'b11111111;
DRAM[9610] = 8'b11111111;
DRAM[9611] = 8'b11111111;
DRAM[9612] = 8'b11111111;
DRAM[9613] = 8'b11111111;
DRAM[9614] = 8'b11111111;
DRAM[9615] = 8'b11111111;
DRAM[9616] = 8'b11111111;
DRAM[9617] = 8'b11111111;
DRAM[9618] = 8'b11111111;
DRAM[9619] = 8'b11111111;
DRAM[9620] = 8'b11111111;
DRAM[9621] = 8'b11111111;
DRAM[9622] = 8'b11111111;
DRAM[9623] = 8'b11111111;
DRAM[9624] = 8'b11111110;
DRAM[9625] = 8'b11111110;
DRAM[9626] = 8'b11111110;
DRAM[9627] = 8'b11111110;
DRAM[9628] = 8'b11111111;
DRAM[9629] = 8'b11111111;
DRAM[9630] = 8'b11111111;
DRAM[9631] = 8'b11111111;
DRAM[9632] = 8'b11111101;
DRAM[9633] = 8'b11111101;
DRAM[9634] = 8'b11111101;
DRAM[9635] = 8'b11111101;
DRAM[9636] = 8'b11111101;
DRAM[9637] = 8'b11111101;
DRAM[9638] = 8'b11111101;
DRAM[9639] = 8'b11111101;
DRAM[9640] = 8'b11111111;
DRAM[9641] = 8'b11111101;
DRAM[9642] = 8'b11111011;
DRAM[9643] = 8'b11111101;
DRAM[9644] = 8'b11111110;
DRAM[9645] = 8'b11111100;
DRAM[9646] = 8'b11111011;
DRAM[9647] = 8'b11111101;
DRAM[9648] = 8'b11111011;
DRAM[9649] = 8'b11111111;
DRAM[9650] = 8'b11101011;
DRAM[9651] = 8'b11100010;
DRAM[9652] = 8'b11010001;
DRAM[9653] = 8'b11000000;
DRAM[9654] = 8'b11010011;
DRAM[9655] = 8'b11001001;
DRAM[9656] = 8'b10100000;
DRAM[9657] = 8'b10110011;
DRAM[9658] = 8'b11011000;
DRAM[9659] = 8'b11110010;
DRAM[9660] = 8'b11011010;
DRAM[9661] = 8'b10100011;
DRAM[9662] = 8'b1111111;
DRAM[9663] = 8'b1111100;
DRAM[9664] = 8'b10100000;
DRAM[9665] = 8'b10010001;
DRAM[9666] = 8'b10000010;
DRAM[9667] = 8'b1110011;
DRAM[9668] = 8'b1101011;
DRAM[9669] = 8'b1110010;
DRAM[9670] = 8'b1110000;
DRAM[9671] = 8'b1011101;
DRAM[9672] = 8'b1100100;
DRAM[9673] = 8'b1100011;
DRAM[9674] = 8'b1100010;
DRAM[9675] = 8'b1100010;
DRAM[9676] = 8'b1100011;
DRAM[9677] = 8'b1100011;
DRAM[9678] = 8'b1100000;
DRAM[9679] = 8'b1011110;
DRAM[9680] = 8'b1011111;
DRAM[9681] = 8'b1011110;
DRAM[9682] = 8'b1011110;
DRAM[9683] = 8'b1011101;
DRAM[9684] = 8'b1011100;
DRAM[9685] = 8'b1011011;
DRAM[9686] = 8'b1011011;
DRAM[9687] = 8'b1011011;
DRAM[9688] = 8'b1011011;
DRAM[9689] = 8'b1011010;
DRAM[9690] = 8'b1011010;
DRAM[9691] = 8'b1011001;
DRAM[9692] = 8'b1011000;
DRAM[9693] = 8'b1010111;
DRAM[9694] = 8'b1010111;
DRAM[9695] = 8'b1010111;
DRAM[9696] = 8'b1010100;
DRAM[9697] = 8'b1010100;
DRAM[9698] = 8'b1010100;
DRAM[9699] = 8'b1010100;
DRAM[9700] = 8'b1010100;
DRAM[9701] = 8'b1010100;
DRAM[9702] = 8'b1010100;
DRAM[9703] = 8'b1010100;
DRAM[9704] = 8'b1010001;
DRAM[9705] = 8'b1010010;
DRAM[9706] = 8'b1010010;
DRAM[9707] = 8'b1010011;
DRAM[9708] = 8'b1010011;
DRAM[9709] = 8'b1010010;
DRAM[9710] = 8'b1010010;
DRAM[9711] = 8'b1010001;
DRAM[9712] = 8'b1010001;
DRAM[9713] = 8'b1010000;
DRAM[9714] = 8'b1010000;
DRAM[9715] = 8'b1010000;
DRAM[9716] = 8'b1001111;
DRAM[9717] = 8'b1001111;
DRAM[9718] = 8'b1001111;
DRAM[9719] = 8'b1001111;
DRAM[9720] = 8'b1001111;
DRAM[9721] = 8'b1001110;
DRAM[9722] = 8'b1001110;
DRAM[9723] = 8'b1001110;
DRAM[9724] = 8'b1001101;
DRAM[9725] = 8'b1001101;
DRAM[9726] = 8'b1001101;
DRAM[9727] = 8'b1001101;
DRAM[9728] = 8'b1100011;
DRAM[9729] = 8'b1100100;
DRAM[9730] = 8'b1100101;
DRAM[9731] = 8'b1100110;
DRAM[9732] = 8'b1100110;
DRAM[9733] = 8'b1100110;
DRAM[9734] = 8'b1100101;
DRAM[9735] = 8'b1100101;
DRAM[9736] = 8'b1101000;
DRAM[9737] = 8'b1101000;
DRAM[9738] = 8'b1101000;
DRAM[9739] = 8'b1101001;
DRAM[9740] = 8'b1101001;
DRAM[9741] = 8'b1101010;
DRAM[9742] = 8'b1101010;
DRAM[9743] = 8'b1101010;
DRAM[9744] = 8'b1101011;
DRAM[9745] = 8'b1101011;
DRAM[9746] = 8'b1101100;
DRAM[9747] = 8'b1101101;
DRAM[9748] = 8'b1101101;
DRAM[9749] = 8'b1101110;
DRAM[9750] = 8'b1101111;
DRAM[9751] = 8'b1101111;
DRAM[9752] = 8'b1101111;
DRAM[9753] = 8'b1101111;
DRAM[9754] = 8'b1110000;
DRAM[9755] = 8'b1110000;
DRAM[9756] = 8'b1110000;
DRAM[9757] = 8'b1110001;
DRAM[9758] = 8'b1110001;
DRAM[9759] = 8'b1110001;
DRAM[9760] = 8'b1110010;
DRAM[9761] = 8'b1110010;
DRAM[9762] = 8'b1110010;
DRAM[9763] = 8'b1110011;
DRAM[9764] = 8'b1110011;
DRAM[9765] = 8'b1110100;
DRAM[9766] = 8'b1110100;
DRAM[9767] = 8'b1110100;
DRAM[9768] = 8'b1110011;
DRAM[9769] = 8'b1110100;
DRAM[9770] = 8'b1110101;
DRAM[9771] = 8'b1110110;
DRAM[9772] = 8'b1110111;
DRAM[9773] = 8'b1111000;
DRAM[9774] = 8'b1111000;
DRAM[9775] = 8'b1110111;
DRAM[9776] = 8'b1111001;
DRAM[9777] = 8'b1111010;
DRAM[9778] = 8'b1111010;
DRAM[9779] = 8'b1111011;
DRAM[9780] = 8'b1111100;
DRAM[9781] = 8'b1111100;
DRAM[9782] = 8'b1111011;
DRAM[9783] = 8'b1111011;
DRAM[9784] = 8'b1111010;
DRAM[9785] = 8'b1111011;
DRAM[9786] = 8'b1111011;
DRAM[9787] = 8'b1111100;
DRAM[9788] = 8'b1111100;
DRAM[9789] = 8'b1111011;
DRAM[9790] = 8'b1111011;
DRAM[9791] = 8'b1111010;
DRAM[9792] = 8'b1111100;
DRAM[9793] = 8'b1111100;
DRAM[9794] = 8'b1111100;
DRAM[9795] = 8'b1111100;
DRAM[9796] = 8'b1111100;
DRAM[9797] = 8'b1111100;
DRAM[9798] = 8'b1111100;
DRAM[9799] = 8'b1111100;
DRAM[9800] = 8'b1111010;
DRAM[9801] = 8'b1111010;
DRAM[9802] = 8'b1111011;
DRAM[9803] = 8'b1111011;
DRAM[9804] = 8'b1111011;
DRAM[9805] = 8'b1111100;
DRAM[9806] = 8'b1111100;
DRAM[9807] = 8'b1111100;
DRAM[9808] = 8'b1111100;
DRAM[9809] = 8'b1111111;
DRAM[9810] = 8'b10000000;
DRAM[9811] = 8'b10000000;
DRAM[9812] = 8'b10000000;
DRAM[9813] = 8'b10000101;
DRAM[9814] = 8'b10001111;
DRAM[9815] = 8'b10010111;
DRAM[9816] = 8'b11000011;
DRAM[9817] = 8'b11000010;
DRAM[9818] = 8'b11011001;
DRAM[9819] = 8'b11110010;
DRAM[9820] = 8'b11101010;
DRAM[9821] = 8'b11111111;
DRAM[9822] = 8'b11111111;
DRAM[9823] = 8'b11111010;
DRAM[9824] = 8'b11111111;
DRAM[9825] = 8'b11111111;
DRAM[9826] = 8'b11111111;
DRAM[9827] = 8'b11111111;
DRAM[9828] = 8'b11111111;
DRAM[9829] = 8'b11111111;
DRAM[9830] = 8'b11111111;
DRAM[9831] = 8'b11111111;
DRAM[9832] = 8'b11111110;
DRAM[9833] = 8'b11111110;
DRAM[9834] = 8'b11111110;
DRAM[9835] = 8'b11111110;
DRAM[9836] = 8'b11111110;
DRAM[9837] = 8'b11111110;
DRAM[9838] = 8'b11111110;
DRAM[9839] = 8'b11111110;
DRAM[9840] = 8'b11111110;
DRAM[9841] = 8'b11111110;
DRAM[9842] = 8'b11111110;
DRAM[9843] = 8'b11111101;
DRAM[9844] = 8'b11111101;
DRAM[9845] = 8'b11111101;
DRAM[9846] = 8'b11111101;
DRAM[9847] = 8'b11111101;
DRAM[9848] = 8'b11111110;
DRAM[9849] = 8'b11111110;
DRAM[9850] = 8'b11111110;
DRAM[9851] = 8'b11111111;
DRAM[9852] = 8'b11111111;
DRAM[9853] = 8'b11111111;
DRAM[9854] = 8'b11111111;
DRAM[9855] = 8'b11111111;
DRAM[9856] = 8'b11111111;
DRAM[9857] = 8'b11111111;
DRAM[9858] = 8'b11111111;
DRAM[9859] = 8'b11111111;
DRAM[9860] = 8'b11111111;
DRAM[9861] = 8'b11111111;
DRAM[9862] = 8'b11111111;
DRAM[9863] = 8'b11111111;
DRAM[9864] = 8'b11111111;
DRAM[9865] = 8'b11111111;
DRAM[9866] = 8'b11111111;
DRAM[9867] = 8'b11111111;
DRAM[9868] = 8'b11111111;
DRAM[9869] = 8'b11111111;
DRAM[9870] = 8'b11111111;
DRAM[9871] = 8'b11111111;
DRAM[9872] = 8'b11111111;
DRAM[9873] = 8'b11111111;
DRAM[9874] = 8'b11111111;
DRAM[9875] = 8'b11111111;
DRAM[9876] = 8'b11111111;
DRAM[9877] = 8'b11111111;
DRAM[9878] = 8'b11111111;
DRAM[9879] = 8'b11111111;
DRAM[9880] = 8'b11111110;
DRAM[9881] = 8'b11111110;
DRAM[9882] = 8'b11111110;
DRAM[9883] = 8'b11111111;
DRAM[9884] = 8'b11111111;
DRAM[9885] = 8'b11111111;
DRAM[9886] = 8'b11111111;
DRAM[9887] = 8'b11111111;
DRAM[9888] = 8'b11111101;
DRAM[9889] = 8'b11111101;
DRAM[9890] = 8'b11111101;
DRAM[9891] = 8'b11111101;
DRAM[9892] = 8'b11111101;
DRAM[9893] = 8'b11111101;
DRAM[9894] = 8'b11111101;
DRAM[9895] = 8'b11111101;
DRAM[9896] = 8'b11111111;
DRAM[9897] = 8'b11111010;
DRAM[9898] = 8'b11111001;
DRAM[9899] = 8'b11111101;
DRAM[9900] = 8'b11111110;
DRAM[9901] = 8'b11111011;
DRAM[9902] = 8'b11111001;
DRAM[9903] = 8'b11111011;
DRAM[9904] = 8'b11111011;
DRAM[9905] = 8'b11111111;
DRAM[9906] = 8'b11101100;
DRAM[9907] = 8'b11111100;
DRAM[9908] = 8'b11111111;
DRAM[9909] = 8'b11111001;
DRAM[9910] = 8'b11111100;
DRAM[9911] = 8'b11100001;
DRAM[9912] = 8'b11110010;
DRAM[9913] = 8'b11111000;
DRAM[9914] = 8'b11111111;
DRAM[9915] = 8'b11110100;
DRAM[9916] = 8'b11010000;
DRAM[9917] = 8'b10101100;
DRAM[9918] = 8'b10100111;
DRAM[9919] = 8'b10110111;
DRAM[9920] = 8'b10111010;
DRAM[9921] = 8'b10001100;
DRAM[9922] = 8'b1110011;
DRAM[9923] = 8'b1111001;
DRAM[9924] = 8'b1111001;
DRAM[9925] = 8'b1110001;
DRAM[9926] = 8'b1101011;
DRAM[9927] = 8'b1100111;
DRAM[9928] = 8'b1100101;
DRAM[9929] = 8'b1100100;
DRAM[9930] = 8'b1100100;
DRAM[9931] = 8'b1100101;
DRAM[9932] = 8'b1100101;
DRAM[9933] = 8'b1100100;
DRAM[9934] = 8'b1100001;
DRAM[9935] = 8'b1011111;
DRAM[9936] = 8'b1011111;
DRAM[9937] = 8'b1011111;
DRAM[9938] = 8'b1011110;
DRAM[9939] = 8'b1011101;
DRAM[9940] = 8'b1011100;
DRAM[9941] = 8'b1011100;
DRAM[9942] = 8'b1011011;
DRAM[9943] = 8'b1011011;
DRAM[9944] = 8'b1011011;
DRAM[9945] = 8'b1011011;
DRAM[9946] = 8'b1011010;
DRAM[9947] = 8'b1011001;
DRAM[9948] = 8'b1011000;
DRAM[9949] = 8'b1011000;
DRAM[9950] = 8'b1010111;
DRAM[9951] = 8'b1010111;
DRAM[9952] = 8'b1010100;
DRAM[9953] = 8'b1010100;
DRAM[9954] = 8'b1010100;
DRAM[9955] = 8'b1010100;
DRAM[9956] = 8'b1010100;
DRAM[9957] = 8'b1010100;
DRAM[9958] = 8'b1010100;
DRAM[9959] = 8'b1010100;
DRAM[9960] = 8'b1010001;
DRAM[9961] = 8'b1010010;
DRAM[9962] = 8'b1010010;
DRAM[9963] = 8'b1010011;
DRAM[9964] = 8'b1010011;
DRAM[9965] = 8'b1010010;
DRAM[9966] = 8'b1010010;
DRAM[9967] = 8'b1010001;
DRAM[9968] = 8'b1010001;
DRAM[9969] = 8'b1010001;
DRAM[9970] = 8'b1010000;
DRAM[9971] = 8'b1010000;
DRAM[9972] = 8'b1010000;
DRAM[9973] = 8'b1001111;
DRAM[9974] = 8'b1001111;
DRAM[9975] = 8'b1001111;
DRAM[9976] = 8'b1001111;
DRAM[9977] = 8'b1001111;
DRAM[9978] = 8'b1001110;
DRAM[9979] = 8'b1001110;
DRAM[9980] = 8'b1001110;
DRAM[9981] = 8'b1001101;
DRAM[9982] = 8'b1001101;
DRAM[9983] = 8'b1001101;
DRAM[9984] = 8'b1100100;
DRAM[9985] = 8'b1100100;
DRAM[9986] = 8'b1100101;
DRAM[9987] = 8'b1100110;
DRAM[9988] = 8'b1100110;
DRAM[9989] = 8'b1100110;
DRAM[9990] = 8'b1100101;
DRAM[9991] = 8'b1100101;
DRAM[9992] = 8'b1101000;
DRAM[9993] = 8'b1101000;
DRAM[9994] = 8'b1101000;
DRAM[9995] = 8'b1101001;
DRAM[9996] = 8'b1101001;
DRAM[9997] = 8'b1101010;
DRAM[9998] = 8'b1101010;
DRAM[9999] = 8'b1101010;
DRAM[10000] = 8'b1101011;
DRAM[10001] = 8'b1101011;
DRAM[10002] = 8'b1101100;
DRAM[10003] = 8'b1101101;
DRAM[10004] = 8'b1101101;
DRAM[10005] = 8'b1101110;
DRAM[10006] = 8'b1101111;
DRAM[10007] = 8'b1101111;
DRAM[10008] = 8'b1101111;
DRAM[10009] = 8'b1101111;
DRAM[10010] = 8'b1101111;
DRAM[10011] = 8'b1110000;
DRAM[10012] = 8'b1110000;
DRAM[10013] = 8'b1110001;
DRAM[10014] = 8'b1110001;
DRAM[10015] = 8'b1110001;
DRAM[10016] = 8'b1110010;
DRAM[10017] = 8'b1110010;
DRAM[10018] = 8'b1110010;
DRAM[10019] = 8'b1110011;
DRAM[10020] = 8'b1110011;
DRAM[10021] = 8'b1110100;
DRAM[10022] = 8'b1110100;
DRAM[10023] = 8'b1110100;
DRAM[10024] = 8'b1110011;
DRAM[10025] = 8'b1110100;
DRAM[10026] = 8'b1110101;
DRAM[10027] = 8'b1110110;
DRAM[10028] = 8'b1110111;
DRAM[10029] = 8'b1111000;
DRAM[10030] = 8'b1111000;
DRAM[10031] = 8'b1111000;
DRAM[10032] = 8'b1111001;
DRAM[10033] = 8'b1111010;
DRAM[10034] = 8'b1111011;
DRAM[10035] = 8'b1111100;
DRAM[10036] = 8'b1111100;
DRAM[10037] = 8'b1111100;
DRAM[10038] = 8'b1111100;
DRAM[10039] = 8'b1111011;
DRAM[10040] = 8'b1111010;
DRAM[10041] = 8'b1111011;
DRAM[10042] = 8'b1111011;
DRAM[10043] = 8'b1111100;
DRAM[10044] = 8'b1111100;
DRAM[10045] = 8'b1111011;
DRAM[10046] = 8'b1111011;
DRAM[10047] = 8'b1111010;
DRAM[10048] = 8'b1111100;
DRAM[10049] = 8'b1111100;
DRAM[10050] = 8'b1111100;
DRAM[10051] = 8'b1111100;
DRAM[10052] = 8'b1111100;
DRAM[10053] = 8'b1111100;
DRAM[10054] = 8'b1111100;
DRAM[10055] = 8'b1111100;
DRAM[10056] = 8'b1111100;
DRAM[10057] = 8'b1111100;
DRAM[10058] = 8'b1111100;
DRAM[10059] = 8'b1111101;
DRAM[10060] = 8'b1111101;
DRAM[10061] = 8'b1111110;
DRAM[10062] = 8'b1111110;
DRAM[10063] = 8'b1111111;
DRAM[10064] = 8'b10000010;
DRAM[10065] = 8'b10000011;
DRAM[10066] = 8'b10000011;
DRAM[10067] = 8'b10000000;
DRAM[10068] = 8'b1111111;
DRAM[10069] = 8'b10000101;
DRAM[10070] = 8'b10001111;
DRAM[10071] = 8'b10011000;
DRAM[10072] = 8'b11001111;
DRAM[10073] = 8'b11110011;
DRAM[10074] = 8'b11101110;
DRAM[10075] = 8'b11111001;
DRAM[10076] = 8'b11111110;
DRAM[10077] = 8'b11111111;
DRAM[10078] = 8'b11101111;
DRAM[10079] = 8'b11111111;
DRAM[10080] = 8'b11111100;
DRAM[10081] = 8'b11111011;
DRAM[10082] = 8'b11111001;
DRAM[10083] = 8'b11111000;
DRAM[10084] = 8'b11111001;
DRAM[10085] = 8'b11111011;
DRAM[10086] = 8'b11111101;
DRAM[10087] = 8'b11111111;
DRAM[10088] = 8'b11111111;
DRAM[10089] = 8'b11111111;
DRAM[10090] = 8'b11111111;
DRAM[10091] = 8'b11111111;
DRAM[10092] = 8'b11111111;
DRAM[10093] = 8'b11111111;
DRAM[10094] = 8'b11111111;
DRAM[10095] = 8'b11111111;
DRAM[10096] = 8'b11111101;
DRAM[10097] = 8'b11111101;
DRAM[10098] = 8'b11111101;
DRAM[10099] = 8'b11111101;
DRAM[10100] = 8'b11111101;
DRAM[10101] = 8'b11111101;
DRAM[10102] = 8'b11111101;
DRAM[10103] = 8'b11111101;
DRAM[10104] = 8'b11111110;
DRAM[10105] = 8'b11111110;
DRAM[10106] = 8'b11111110;
DRAM[10107] = 8'b11111111;
DRAM[10108] = 8'b11111111;
DRAM[10109] = 8'b11111111;
DRAM[10110] = 8'b11111111;
DRAM[10111] = 8'b11111111;
DRAM[10112] = 8'b11111111;
DRAM[10113] = 8'b11111111;
DRAM[10114] = 8'b11111111;
DRAM[10115] = 8'b11111111;
DRAM[10116] = 8'b11111111;
DRAM[10117] = 8'b11111111;
DRAM[10118] = 8'b11111111;
DRAM[10119] = 8'b11111111;
DRAM[10120] = 8'b11111111;
DRAM[10121] = 8'b11111111;
DRAM[10122] = 8'b11111111;
DRAM[10123] = 8'b11111111;
DRAM[10124] = 8'b11111111;
DRAM[10125] = 8'b11111111;
DRAM[10126] = 8'b11111111;
DRAM[10127] = 8'b11111111;
DRAM[10128] = 8'b11111111;
DRAM[10129] = 8'b11111111;
DRAM[10130] = 8'b11111111;
DRAM[10131] = 8'b11111111;
DRAM[10132] = 8'b11111111;
DRAM[10133] = 8'b11111111;
DRAM[10134] = 8'b11111111;
DRAM[10135] = 8'b11111111;
DRAM[10136] = 8'b11111110;
DRAM[10137] = 8'b11111110;
DRAM[10138] = 8'b11111110;
DRAM[10139] = 8'b11111111;
DRAM[10140] = 8'b11111111;
DRAM[10141] = 8'b11111111;
DRAM[10142] = 8'b11111111;
DRAM[10143] = 8'b11111111;
DRAM[10144] = 8'b11111110;
DRAM[10145] = 8'b11111110;
DRAM[10146] = 8'b11111110;
DRAM[10147] = 8'b11111110;
DRAM[10148] = 8'b11111110;
DRAM[10149] = 8'b11111110;
DRAM[10150] = 8'b11111110;
DRAM[10151] = 8'b11111110;
DRAM[10152] = 8'b11111111;
DRAM[10153] = 8'b11111100;
DRAM[10154] = 8'b11111100;
DRAM[10155] = 8'b11111111;
DRAM[10156] = 8'b11111111;
DRAM[10157] = 8'b11111011;
DRAM[10158] = 8'b11111001;
DRAM[10159] = 8'b11111100;
DRAM[10160] = 8'b11111111;
DRAM[10161] = 8'b11110010;
DRAM[10162] = 8'b11111111;
DRAM[10163] = 8'b11110110;
DRAM[10164] = 8'b11110001;
DRAM[10165] = 8'b11111000;
DRAM[10166] = 8'b11101011;
DRAM[10167] = 8'b11111111;
DRAM[10168] = 8'b11110111;
DRAM[10169] = 8'b11110111;
DRAM[10170] = 8'b11110110;
DRAM[10171] = 8'b11110100;
DRAM[10172] = 8'b11101111;
DRAM[10173] = 8'b11100111;
DRAM[10174] = 8'b11011110;
DRAM[10175] = 8'b11010111;
DRAM[10176] = 8'b10101100;
DRAM[10177] = 8'b1111101;
DRAM[10178] = 8'b1111010;
DRAM[10179] = 8'b10011111;
DRAM[10180] = 8'b10011101;
DRAM[10181] = 8'b1110110;
DRAM[10182] = 8'b1100011;
DRAM[10183] = 8'b1101011;
DRAM[10184] = 8'b1100111;
DRAM[10185] = 8'b1100110;
DRAM[10186] = 8'b1100110;
DRAM[10187] = 8'b1100110;
DRAM[10188] = 8'b1100111;
DRAM[10189] = 8'b1100110;
DRAM[10190] = 8'b1100011;
DRAM[10191] = 8'b1100000;
DRAM[10192] = 8'b1011111;
DRAM[10193] = 8'b1011111;
DRAM[10194] = 8'b1011110;
DRAM[10195] = 8'b1011101;
DRAM[10196] = 8'b1011101;
DRAM[10197] = 8'b1011100;
DRAM[10198] = 8'b1011011;
DRAM[10199] = 8'b1011011;
DRAM[10200] = 8'b1011011;
DRAM[10201] = 8'b1011011;
DRAM[10202] = 8'b1011010;
DRAM[10203] = 8'b1011001;
DRAM[10204] = 8'b1011001;
DRAM[10205] = 8'b1011000;
DRAM[10206] = 8'b1010111;
DRAM[10207] = 8'b1010111;
DRAM[10208] = 8'b1010100;
DRAM[10209] = 8'b1010100;
DRAM[10210] = 8'b1010100;
DRAM[10211] = 8'b1010100;
DRAM[10212] = 8'b1010100;
DRAM[10213] = 8'b1010100;
DRAM[10214] = 8'b1010100;
DRAM[10215] = 8'b1010100;
DRAM[10216] = 8'b1010001;
DRAM[10217] = 8'b1010010;
DRAM[10218] = 8'b1010010;
DRAM[10219] = 8'b1010011;
DRAM[10220] = 8'b1010011;
DRAM[10221] = 8'b1010010;
DRAM[10222] = 8'b1010010;
DRAM[10223] = 8'b1010001;
DRAM[10224] = 8'b1010001;
DRAM[10225] = 8'b1010001;
DRAM[10226] = 8'b1010001;
DRAM[10227] = 8'b1010000;
DRAM[10228] = 8'b1010000;
DRAM[10229] = 8'b1001111;
DRAM[10230] = 8'b1001111;
DRAM[10231] = 8'b1001111;
DRAM[10232] = 8'b1001111;
DRAM[10233] = 8'b1001111;
DRAM[10234] = 8'b1001111;
DRAM[10235] = 8'b1001110;
DRAM[10236] = 8'b1001110;
DRAM[10237] = 8'b1001101;
DRAM[10238] = 8'b1001101;
DRAM[10239] = 8'b1001101;
DRAM[10240] = 8'b1100100;
DRAM[10241] = 8'b1100100;
DRAM[10242] = 8'b1100101;
DRAM[10243] = 8'b1100110;
DRAM[10244] = 8'b1100110;
DRAM[10245] = 8'b1100111;
DRAM[10246] = 8'b1101000;
DRAM[10247] = 8'b1101000;
DRAM[10248] = 8'b1100110;
DRAM[10249] = 8'b1100110;
DRAM[10250] = 8'b1100111;
DRAM[10251] = 8'b1101000;
DRAM[10252] = 8'b1101000;
DRAM[10253] = 8'b1101001;
DRAM[10254] = 8'b1101010;
DRAM[10255] = 8'b1101010;
DRAM[10256] = 8'b1101010;
DRAM[10257] = 8'b1101010;
DRAM[10258] = 8'b1101011;
DRAM[10259] = 8'b1101100;
DRAM[10260] = 8'b1101100;
DRAM[10261] = 8'b1101101;
DRAM[10262] = 8'b1101110;
DRAM[10263] = 8'b1101110;
DRAM[10264] = 8'b1101011;
DRAM[10265] = 8'b1101101;
DRAM[10266] = 8'b1101110;
DRAM[10267] = 8'b1110000;
DRAM[10268] = 8'b1110001;
DRAM[10269] = 8'b1110001;
DRAM[10270] = 8'b1110000;
DRAM[10271] = 8'b1101111;
DRAM[10272] = 8'b1110011;
DRAM[10273] = 8'b1110011;
DRAM[10274] = 8'b1110011;
DRAM[10275] = 8'b1110100;
DRAM[10276] = 8'b1110100;
DRAM[10277] = 8'b1110101;
DRAM[10278] = 8'b1110101;
DRAM[10279] = 8'b1110101;
DRAM[10280] = 8'b1110100;
DRAM[10281] = 8'b1110100;
DRAM[10282] = 8'b1110101;
DRAM[10283] = 8'b1110110;
DRAM[10284] = 8'b1110110;
DRAM[10285] = 8'b1110111;
DRAM[10286] = 8'b1111000;
DRAM[10287] = 8'b1111000;
DRAM[10288] = 8'b1111001;
DRAM[10289] = 8'b1111001;
DRAM[10290] = 8'b1111000;
DRAM[10291] = 8'b1111010;
DRAM[10292] = 8'b1111100;
DRAM[10293] = 8'b1111100;
DRAM[10294] = 8'b1111011;
DRAM[10295] = 8'b1111001;
DRAM[10296] = 8'b1111011;
DRAM[10297] = 8'b1111100;
DRAM[10298] = 8'b1111100;
DRAM[10299] = 8'b1111100;
DRAM[10300] = 8'b1111011;
DRAM[10301] = 8'b1111010;
DRAM[10302] = 8'b1111001;
DRAM[10303] = 8'b1111001;
DRAM[10304] = 8'b1111010;
DRAM[10305] = 8'b1111100;
DRAM[10306] = 8'b10000000;
DRAM[10307] = 8'b10000001;
DRAM[10308] = 8'b1111101;
DRAM[10309] = 8'b1111001;
DRAM[10310] = 8'b1111011;
DRAM[10311] = 8'b1111111;
DRAM[10312] = 8'b1111100;
DRAM[10313] = 8'b10000011;
DRAM[10314] = 8'b1111011;
DRAM[10315] = 8'b1110011;
DRAM[10316] = 8'b1111100;
DRAM[10317] = 8'b10000010;
DRAM[10318] = 8'b10000001;
DRAM[10319] = 8'b10000011;
DRAM[10320] = 8'b10000101;
DRAM[10321] = 8'b10001001;
DRAM[10322] = 8'b10001001;
DRAM[10323] = 8'b10000110;
DRAM[10324] = 8'b10001110;
DRAM[10325] = 8'b10100110;
DRAM[10326] = 8'b11000100;
DRAM[10327] = 8'b11010111;
DRAM[10328] = 8'b11101100;
DRAM[10329] = 8'b11110000;
DRAM[10330] = 8'b11110110;
DRAM[10331] = 8'b11111011;
DRAM[10332] = 8'b11111110;
DRAM[10333] = 8'b11111111;
DRAM[10334] = 8'b11111110;
DRAM[10335] = 8'b11111101;
DRAM[10336] = 8'b11111111;
DRAM[10337] = 8'b11111111;
DRAM[10338] = 8'b11111111;
DRAM[10339] = 8'b11111111;
DRAM[10340] = 8'b11111111;
DRAM[10341] = 8'b11111111;
DRAM[10342] = 8'b11111111;
DRAM[10343] = 8'b11111111;
DRAM[10344] = 8'b11111110;
DRAM[10345] = 8'b11111110;
DRAM[10346] = 8'b11111110;
DRAM[10347] = 8'b11111110;
DRAM[10348] = 8'b11111110;
DRAM[10349] = 8'b11111110;
DRAM[10350] = 8'b11111110;
DRAM[10351] = 8'b11111110;
DRAM[10352] = 8'b11111110;
DRAM[10353] = 8'b11111110;
DRAM[10354] = 8'b11111110;
DRAM[10355] = 8'b11111110;
DRAM[10356] = 8'b11111110;
DRAM[10357] = 8'b11111110;
DRAM[10358] = 8'b11111110;
DRAM[10359] = 8'b11111110;
DRAM[10360] = 8'b11111110;
DRAM[10361] = 8'b11111110;
DRAM[10362] = 8'b11111110;
DRAM[10363] = 8'b11111111;
DRAM[10364] = 8'b11111111;
DRAM[10365] = 8'b11111111;
DRAM[10366] = 8'b11111111;
DRAM[10367] = 8'b11111111;
DRAM[10368] = 8'b11111111;
DRAM[10369] = 8'b11111111;
DRAM[10370] = 8'b11111111;
DRAM[10371] = 8'b11111111;
DRAM[10372] = 8'b11111111;
DRAM[10373] = 8'b11111111;
DRAM[10374] = 8'b11111111;
DRAM[10375] = 8'b11111111;
DRAM[10376] = 8'b11111111;
DRAM[10377] = 8'b11111111;
DRAM[10378] = 8'b11111111;
DRAM[10379] = 8'b11111111;
DRAM[10380] = 8'b11111111;
DRAM[10381] = 8'b11111111;
DRAM[10382] = 8'b11111111;
DRAM[10383] = 8'b11111111;
DRAM[10384] = 8'b11111101;
DRAM[10385] = 8'b11111101;
DRAM[10386] = 8'b11111101;
DRAM[10387] = 8'b11111110;
DRAM[10388] = 8'b11111110;
DRAM[10389] = 8'b11111111;
DRAM[10390] = 8'b11111111;
DRAM[10391] = 8'b11111111;
DRAM[10392] = 8'b11111110;
DRAM[10393] = 8'b11111110;
DRAM[10394] = 8'b11111110;
DRAM[10395] = 8'b11111111;
DRAM[10396] = 8'b11111111;
DRAM[10397] = 8'b11111111;
DRAM[10398] = 8'b11111111;
DRAM[10399] = 8'b11111111;
DRAM[10400] = 8'b11111110;
DRAM[10401] = 8'b11111110;
DRAM[10402] = 8'b11111110;
DRAM[10403] = 8'b11111110;
DRAM[10404] = 8'b11111110;
DRAM[10405] = 8'b11111110;
DRAM[10406] = 8'b11111110;
DRAM[10407] = 8'b11111110;
DRAM[10408] = 8'b11111101;
DRAM[10409] = 8'b11111101;
DRAM[10410] = 8'b11111101;
DRAM[10411] = 8'b11111110;
DRAM[10412] = 8'b11111110;
DRAM[10413] = 8'b11111111;
DRAM[10414] = 8'b11111111;
DRAM[10415] = 8'b11111111;
DRAM[10416] = 8'b11111100;
DRAM[10417] = 8'b11111100;
DRAM[10418] = 8'b11111100;
DRAM[10419] = 8'b11111100;
DRAM[10420] = 8'b11111100;
DRAM[10421] = 8'b11111100;
DRAM[10422] = 8'b11111100;
DRAM[10423] = 8'b11111100;
DRAM[10424] = 8'b11111010;
DRAM[10425] = 8'b11111111;
DRAM[10426] = 8'b11111101;
DRAM[10427] = 8'b11110111;
DRAM[10428] = 8'b11111001;
DRAM[10429] = 8'b11111011;
DRAM[10430] = 8'b11101111;
DRAM[10431] = 8'b11011100;
DRAM[10432] = 8'b10100001;
DRAM[10433] = 8'b10010100;
DRAM[10434] = 8'b10110100;
DRAM[10435] = 8'b11000101;
DRAM[10436] = 8'b10010101;
DRAM[10437] = 8'b1101111;
DRAM[10438] = 8'b1110101;
DRAM[10439] = 8'b1111011;
DRAM[10440] = 8'b1111010;
DRAM[10441] = 8'b1110011;
DRAM[10442] = 8'b1101101;
DRAM[10443] = 8'b1101100;
DRAM[10444] = 8'b1101111;
DRAM[10445] = 8'b1110001;
DRAM[10446] = 8'b1101101;
DRAM[10447] = 8'b1101000;
DRAM[10448] = 8'b1100010;
DRAM[10449] = 8'b1100010;
DRAM[10450] = 8'b1100001;
DRAM[10451] = 8'b1011110;
DRAM[10452] = 8'b1011011;
DRAM[10453] = 8'b1011010;
DRAM[10454] = 8'b1011010;
DRAM[10455] = 8'b1011011;
DRAM[10456] = 8'b1011010;
DRAM[10457] = 8'b1011010;
DRAM[10458] = 8'b1011001;
DRAM[10459] = 8'b1011000;
DRAM[10460] = 8'b1011000;
DRAM[10461] = 8'b1010111;
DRAM[10462] = 8'b1010110;
DRAM[10463] = 8'b1010110;
DRAM[10464] = 8'b1010110;
DRAM[10465] = 8'b1010110;
DRAM[10466] = 8'b1010110;
DRAM[10467] = 8'b1010101;
DRAM[10468] = 8'b1010101;
DRAM[10469] = 8'b1010100;
DRAM[10470] = 8'b1010100;
DRAM[10471] = 8'b1010100;
DRAM[10472] = 8'b1010001;
DRAM[10473] = 8'b1010010;
DRAM[10474] = 8'b1010010;
DRAM[10475] = 8'b1010011;
DRAM[10476] = 8'b1010011;
DRAM[10477] = 8'b1010010;
DRAM[10478] = 8'b1010010;
DRAM[10479] = 8'b1010001;
DRAM[10480] = 8'b1010010;
DRAM[10481] = 8'b1010010;
DRAM[10482] = 8'b1010010;
DRAM[10483] = 8'b1010001;
DRAM[10484] = 8'b1010001;
DRAM[10485] = 8'b1010000;
DRAM[10486] = 8'b1010000;
DRAM[10487] = 8'b1010000;
DRAM[10488] = 8'b1010000;
DRAM[10489] = 8'b1010000;
DRAM[10490] = 8'b1010000;
DRAM[10491] = 8'b1010000;
DRAM[10492] = 8'b1010000;
DRAM[10493] = 8'b1010000;
DRAM[10494] = 8'b1010000;
DRAM[10495] = 8'b1010000;
DRAM[10496] = 8'b1100011;
DRAM[10497] = 8'b1100011;
DRAM[10498] = 8'b1100100;
DRAM[10499] = 8'b1100100;
DRAM[10500] = 8'b1100101;
DRAM[10501] = 8'b1100110;
DRAM[10502] = 8'b1100111;
DRAM[10503] = 8'b1100111;
DRAM[10504] = 8'b1100110;
DRAM[10505] = 8'b1100110;
DRAM[10506] = 8'b1100111;
DRAM[10507] = 8'b1101000;
DRAM[10508] = 8'b1101000;
DRAM[10509] = 8'b1101001;
DRAM[10510] = 8'b1101010;
DRAM[10511] = 8'b1101010;
DRAM[10512] = 8'b1101010;
DRAM[10513] = 8'b1101010;
DRAM[10514] = 8'b1101011;
DRAM[10515] = 8'b1101100;
DRAM[10516] = 8'b1101100;
DRAM[10517] = 8'b1101101;
DRAM[10518] = 8'b1101110;
DRAM[10519] = 8'b1101110;
DRAM[10520] = 8'b1101100;
DRAM[10521] = 8'b1101101;
DRAM[10522] = 8'b1101110;
DRAM[10523] = 8'b1110000;
DRAM[10524] = 8'b1110001;
DRAM[10525] = 8'b1110001;
DRAM[10526] = 8'b1110000;
DRAM[10527] = 8'b1110000;
DRAM[10528] = 8'b1110011;
DRAM[10529] = 8'b1110011;
DRAM[10530] = 8'b1110011;
DRAM[10531] = 8'b1110100;
DRAM[10532] = 8'b1110100;
DRAM[10533] = 8'b1110101;
DRAM[10534] = 8'b1110101;
DRAM[10535] = 8'b1110101;
DRAM[10536] = 8'b1110100;
DRAM[10537] = 8'b1110100;
DRAM[10538] = 8'b1110101;
DRAM[10539] = 8'b1110110;
DRAM[10540] = 8'b1110110;
DRAM[10541] = 8'b1110111;
DRAM[10542] = 8'b1111000;
DRAM[10543] = 8'b1111000;
DRAM[10544] = 8'b1111001;
DRAM[10545] = 8'b1111001;
DRAM[10546] = 8'b1111000;
DRAM[10547] = 8'b1111010;
DRAM[10548] = 8'b1111100;
DRAM[10549] = 8'b1111100;
DRAM[10550] = 8'b1111011;
DRAM[10551] = 8'b1111001;
DRAM[10552] = 8'b1111011;
DRAM[10553] = 8'b1111011;
DRAM[10554] = 8'b1111100;
DRAM[10555] = 8'b1111101;
DRAM[10556] = 8'b1111101;
DRAM[10557] = 8'b1111110;
DRAM[10558] = 8'b1111110;
DRAM[10559] = 8'b1111101;
DRAM[10560] = 8'b10000010;
DRAM[10561] = 8'b1111100;
DRAM[10562] = 8'b1110111;
DRAM[10563] = 8'b1111000;
DRAM[10564] = 8'b1111100;
DRAM[10565] = 8'b1111111;
DRAM[10566] = 8'b10000000;
DRAM[10567] = 8'b10000000;
DRAM[10568] = 8'b10001000;
DRAM[10569] = 8'b1111100;
DRAM[10570] = 8'b1110111;
DRAM[10571] = 8'b10001000;
DRAM[10572] = 8'b10010001;
DRAM[10573] = 8'b10000000;
DRAM[10574] = 8'b1111011;
DRAM[10575] = 8'b10010001;
DRAM[10576] = 8'b10100111;
DRAM[10577] = 8'b10101110;
DRAM[10578] = 8'b10110001;
DRAM[10579] = 8'b10101101;
DRAM[10580] = 8'b10110010;
DRAM[10581] = 8'b11001011;
DRAM[10582] = 8'b11101100;
DRAM[10583] = 8'b11111111;
DRAM[10584] = 8'b11110100;
DRAM[10585] = 8'b11110110;
DRAM[10586] = 8'b11111010;
DRAM[10587] = 8'b11111101;
DRAM[10588] = 8'b11111111;
DRAM[10589] = 8'b11111111;
DRAM[10590] = 8'b11111110;
DRAM[10591] = 8'b11111101;
DRAM[10592] = 8'b11111111;
DRAM[10593] = 8'b11111111;
DRAM[10594] = 8'b11111111;
DRAM[10595] = 8'b11111111;
DRAM[10596] = 8'b11111111;
DRAM[10597] = 8'b11111111;
DRAM[10598] = 8'b11111111;
DRAM[10599] = 8'b11111111;
DRAM[10600] = 8'b11111110;
DRAM[10601] = 8'b11111110;
DRAM[10602] = 8'b11111110;
DRAM[10603] = 8'b11111110;
DRAM[10604] = 8'b11111110;
DRAM[10605] = 8'b11111110;
DRAM[10606] = 8'b11111110;
DRAM[10607] = 8'b11111110;
DRAM[10608] = 8'b11111110;
DRAM[10609] = 8'b11111110;
DRAM[10610] = 8'b11111110;
DRAM[10611] = 8'b11111110;
DRAM[10612] = 8'b11111110;
DRAM[10613] = 8'b11111110;
DRAM[10614] = 8'b11111110;
DRAM[10615] = 8'b11111110;
DRAM[10616] = 8'b11111110;
DRAM[10617] = 8'b11111110;
DRAM[10618] = 8'b11111110;
DRAM[10619] = 8'b11111111;
DRAM[10620] = 8'b11111111;
DRAM[10621] = 8'b11111111;
DRAM[10622] = 8'b11111111;
DRAM[10623] = 8'b11111111;
DRAM[10624] = 8'b11111111;
DRAM[10625] = 8'b11111111;
DRAM[10626] = 8'b11111111;
DRAM[10627] = 8'b11111111;
DRAM[10628] = 8'b11111111;
DRAM[10629] = 8'b11111111;
DRAM[10630] = 8'b11111111;
DRAM[10631] = 8'b11111111;
DRAM[10632] = 8'b11111111;
DRAM[10633] = 8'b11111111;
DRAM[10634] = 8'b11111111;
DRAM[10635] = 8'b11111111;
DRAM[10636] = 8'b11111111;
DRAM[10637] = 8'b11111111;
DRAM[10638] = 8'b11111111;
DRAM[10639] = 8'b11111111;
DRAM[10640] = 8'b11111101;
DRAM[10641] = 8'b11111101;
DRAM[10642] = 8'b11111101;
DRAM[10643] = 8'b11111110;
DRAM[10644] = 8'b11111110;
DRAM[10645] = 8'b11111111;
DRAM[10646] = 8'b11111111;
DRAM[10647] = 8'b11111111;
DRAM[10648] = 8'b11111110;
DRAM[10649] = 8'b11111110;
DRAM[10650] = 8'b11111110;
DRAM[10651] = 8'b11111111;
DRAM[10652] = 8'b11111111;
DRAM[10653] = 8'b11111111;
DRAM[10654] = 8'b11111111;
DRAM[10655] = 8'b11111111;
DRAM[10656] = 8'b11111110;
DRAM[10657] = 8'b11111110;
DRAM[10658] = 8'b11111110;
DRAM[10659] = 8'b11111110;
DRAM[10660] = 8'b11111110;
DRAM[10661] = 8'b11111110;
DRAM[10662] = 8'b11111110;
DRAM[10663] = 8'b11111110;
DRAM[10664] = 8'b11111101;
DRAM[10665] = 8'b11111101;
DRAM[10666] = 8'b11111101;
DRAM[10667] = 8'b11111110;
DRAM[10668] = 8'b11111110;
DRAM[10669] = 8'b11111111;
DRAM[10670] = 8'b11111111;
DRAM[10671] = 8'b11111111;
DRAM[10672] = 8'b11111110;
DRAM[10673] = 8'b11111110;
DRAM[10674] = 8'b11111110;
DRAM[10675] = 8'b11111110;
DRAM[10676] = 8'b11111110;
DRAM[10677] = 8'b11111110;
DRAM[10678] = 8'b11111110;
DRAM[10679] = 8'b11111110;
DRAM[10680] = 8'b11111100;
DRAM[10681] = 8'b11111111;
DRAM[10682] = 8'b11111110;
DRAM[10683] = 8'b11111001;
DRAM[10684] = 8'b11111011;
DRAM[10685] = 8'b11111110;
DRAM[10686] = 8'b11110100;
DRAM[10687] = 8'b11100100;
DRAM[10688] = 8'b11000011;
DRAM[10689] = 8'b11000100;
DRAM[10690] = 8'b11011101;
DRAM[10691] = 8'b11010111;
DRAM[10692] = 8'b10100011;
DRAM[10693] = 8'b10001000;
DRAM[10694] = 8'b10010000;
DRAM[10695] = 8'b10001111;
DRAM[10696] = 8'b10001001;
DRAM[10697] = 8'b1111110;
DRAM[10698] = 8'b1110010;
DRAM[10699] = 8'b1101110;
DRAM[10700] = 8'b1101111;
DRAM[10701] = 8'b1101100;
DRAM[10702] = 8'b1100011;
DRAM[10703] = 8'b1011011;
DRAM[10704] = 8'b1100011;
DRAM[10705] = 8'b1100010;
DRAM[10706] = 8'b1100010;
DRAM[10707] = 8'b1100000;
DRAM[10708] = 8'b1011101;
DRAM[10709] = 8'b1011100;
DRAM[10710] = 8'b1011011;
DRAM[10711] = 8'b1011011;
DRAM[10712] = 8'b1011010;
DRAM[10713] = 8'b1011010;
DRAM[10714] = 8'b1011001;
DRAM[10715] = 8'b1011001;
DRAM[10716] = 8'b1011000;
DRAM[10717] = 8'b1010111;
DRAM[10718] = 8'b1010110;
DRAM[10719] = 8'b1010110;
DRAM[10720] = 8'b1010110;
DRAM[10721] = 8'b1010110;
DRAM[10722] = 8'b1010110;
DRAM[10723] = 8'b1010101;
DRAM[10724] = 8'b1010101;
DRAM[10725] = 8'b1010100;
DRAM[10726] = 8'b1010100;
DRAM[10727] = 8'b1010100;
DRAM[10728] = 8'b1010001;
DRAM[10729] = 8'b1010010;
DRAM[10730] = 8'b1010010;
DRAM[10731] = 8'b1010011;
DRAM[10732] = 8'b1010011;
DRAM[10733] = 8'b1010010;
DRAM[10734] = 8'b1010010;
DRAM[10735] = 8'b1010001;
DRAM[10736] = 8'b1010010;
DRAM[10737] = 8'b1010010;
DRAM[10738] = 8'b1010010;
DRAM[10739] = 8'b1010001;
DRAM[10740] = 8'b1010001;
DRAM[10741] = 8'b1010000;
DRAM[10742] = 8'b1010000;
DRAM[10743] = 8'b1010000;
DRAM[10744] = 8'b1001111;
DRAM[10745] = 8'b1001111;
DRAM[10746] = 8'b1001111;
DRAM[10747] = 8'b1001111;
DRAM[10748] = 8'b1001111;
DRAM[10749] = 8'b1001111;
DRAM[10750] = 8'b1001111;
DRAM[10751] = 8'b1001111;
DRAM[10752] = 8'b1100010;
DRAM[10753] = 8'b1100010;
DRAM[10754] = 8'b1100011;
DRAM[10755] = 8'b1100011;
DRAM[10756] = 8'b1100100;
DRAM[10757] = 8'b1100101;
DRAM[10758] = 8'b1100110;
DRAM[10759] = 8'b1100110;
DRAM[10760] = 8'b1100110;
DRAM[10761] = 8'b1100110;
DRAM[10762] = 8'b1100111;
DRAM[10763] = 8'b1101000;
DRAM[10764] = 8'b1101000;
DRAM[10765] = 8'b1101001;
DRAM[10766] = 8'b1101010;
DRAM[10767] = 8'b1101010;
DRAM[10768] = 8'b1101010;
DRAM[10769] = 8'b1101010;
DRAM[10770] = 8'b1101011;
DRAM[10771] = 8'b1101100;
DRAM[10772] = 8'b1101100;
DRAM[10773] = 8'b1101101;
DRAM[10774] = 8'b1101110;
DRAM[10775] = 8'b1101110;
DRAM[10776] = 8'b1101100;
DRAM[10777] = 8'b1101101;
DRAM[10778] = 8'b1101110;
DRAM[10779] = 8'b1101111;
DRAM[10780] = 8'b1110000;
DRAM[10781] = 8'b1110001;
DRAM[10782] = 8'b1110000;
DRAM[10783] = 8'b1110000;
DRAM[10784] = 8'b1110011;
DRAM[10785] = 8'b1110011;
DRAM[10786] = 8'b1110011;
DRAM[10787] = 8'b1110100;
DRAM[10788] = 8'b1110100;
DRAM[10789] = 8'b1110101;
DRAM[10790] = 8'b1110101;
DRAM[10791] = 8'b1110101;
DRAM[10792] = 8'b1110100;
DRAM[10793] = 8'b1110100;
DRAM[10794] = 8'b1110101;
DRAM[10795] = 8'b1110110;
DRAM[10796] = 8'b1110110;
DRAM[10797] = 8'b1110111;
DRAM[10798] = 8'b1111000;
DRAM[10799] = 8'b1111000;
DRAM[10800] = 8'b1111001;
DRAM[10801] = 8'b1111001;
DRAM[10802] = 8'b1111000;
DRAM[10803] = 8'b1111010;
DRAM[10804] = 8'b1111100;
DRAM[10805] = 8'b1111100;
DRAM[10806] = 8'b1111011;
DRAM[10807] = 8'b1111001;
DRAM[10808] = 8'b1111011;
DRAM[10809] = 8'b1111011;
DRAM[10810] = 8'b1111100;
DRAM[10811] = 8'b1111100;
DRAM[10812] = 8'b1111101;
DRAM[10813] = 8'b1111110;
DRAM[10814] = 8'b1111110;
DRAM[10815] = 8'b1111111;
DRAM[10816] = 8'b1110110;
DRAM[10817] = 8'b1111011;
DRAM[10818] = 8'b10000010;
DRAM[10819] = 8'b10000111;
DRAM[10820] = 8'b10001001;
DRAM[10821] = 8'b10000111;
DRAM[10822] = 8'b10000011;
DRAM[10823] = 8'b1111111;
DRAM[10824] = 8'b10000110;
DRAM[10825] = 8'b10001011;
DRAM[10826] = 8'b10001001;
DRAM[10827] = 8'b10001001;
DRAM[10828] = 8'b10010000;
DRAM[10829] = 8'b10001100;
DRAM[10830] = 8'b10000100;
DRAM[10831] = 8'b10000110;
DRAM[10832] = 8'b10001111;
DRAM[10833] = 8'b10110011;
DRAM[10834] = 8'b11011110;
DRAM[10835] = 8'b11110101;
DRAM[10836] = 8'b11111011;
DRAM[10837] = 8'b11111011;
DRAM[10838] = 8'b11111010;
DRAM[10839] = 8'b11111001;
DRAM[10840] = 8'b11111101;
DRAM[10841] = 8'b11111110;
DRAM[10842] = 8'b11111111;
DRAM[10843] = 8'b11111111;
DRAM[10844] = 8'b11111111;
DRAM[10845] = 8'b11111111;
DRAM[10846] = 8'b11111111;
DRAM[10847] = 8'b11111111;
DRAM[10848] = 8'b11111111;
DRAM[10849] = 8'b11111111;
DRAM[10850] = 8'b11111111;
DRAM[10851] = 8'b11111111;
DRAM[10852] = 8'b11111111;
DRAM[10853] = 8'b11111111;
DRAM[10854] = 8'b11111111;
DRAM[10855] = 8'b11111111;
DRAM[10856] = 8'b11111110;
DRAM[10857] = 8'b11111110;
DRAM[10858] = 8'b11111110;
DRAM[10859] = 8'b11111110;
DRAM[10860] = 8'b11111110;
DRAM[10861] = 8'b11111110;
DRAM[10862] = 8'b11111110;
DRAM[10863] = 8'b11111110;
DRAM[10864] = 8'b11111110;
DRAM[10865] = 8'b11111110;
DRAM[10866] = 8'b11111110;
DRAM[10867] = 8'b11111110;
DRAM[10868] = 8'b11111110;
DRAM[10869] = 8'b11111110;
DRAM[10870] = 8'b11111110;
DRAM[10871] = 8'b11111110;
DRAM[10872] = 8'b11111110;
DRAM[10873] = 8'b11111110;
DRAM[10874] = 8'b11111110;
DRAM[10875] = 8'b11111111;
DRAM[10876] = 8'b11111111;
DRAM[10877] = 8'b11111111;
DRAM[10878] = 8'b11111111;
DRAM[10879] = 8'b11111111;
DRAM[10880] = 8'b11111111;
DRAM[10881] = 8'b11111111;
DRAM[10882] = 8'b11111111;
DRAM[10883] = 8'b11111111;
DRAM[10884] = 8'b11111111;
DRAM[10885] = 8'b11111111;
DRAM[10886] = 8'b11111111;
DRAM[10887] = 8'b11111111;
DRAM[10888] = 8'b11111111;
DRAM[10889] = 8'b11111111;
DRAM[10890] = 8'b11111111;
DRAM[10891] = 8'b11111111;
DRAM[10892] = 8'b11111111;
DRAM[10893] = 8'b11111111;
DRAM[10894] = 8'b11111111;
DRAM[10895] = 8'b11111111;
DRAM[10896] = 8'b11111101;
DRAM[10897] = 8'b11111101;
DRAM[10898] = 8'b11111110;
DRAM[10899] = 8'b11111110;
DRAM[10900] = 8'b11111110;
DRAM[10901] = 8'b11111110;
DRAM[10902] = 8'b11111111;
DRAM[10903] = 8'b11111111;
DRAM[10904] = 8'b11111110;
DRAM[10905] = 8'b11111110;
DRAM[10906] = 8'b11111110;
DRAM[10907] = 8'b11111111;
DRAM[10908] = 8'b11111111;
DRAM[10909] = 8'b11111111;
DRAM[10910] = 8'b11111111;
DRAM[10911] = 8'b11111111;
DRAM[10912] = 8'b11111110;
DRAM[10913] = 8'b11111110;
DRAM[10914] = 8'b11111110;
DRAM[10915] = 8'b11111110;
DRAM[10916] = 8'b11111110;
DRAM[10917] = 8'b11111110;
DRAM[10918] = 8'b11111110;
DRAM[10919] = 8'b11111110;
DRAM[10920] = 8'b11111101;
DRAM[10921] = 8'b11111101;
DRAM[10922] = 8'b11111101;
DRAM[10923] = 8'b11111110;
DRAM[10924] = 8'b11111110;
DRAM[10925] = 8'b11111111;
DRAM[10926] = 8'b11111111;
DRAM[10927] = 8'b11111111;
DRAM[10928] = 8'b11111111;
DRAM[10929] = 8'b11111111;
DRAM[10930] = 8'b11111111;
DRAM[10931] = 8'b11111111;
DRAM[10932] = 8'b11111111;
DRAM[10933] = 8'b11111111;
DRAM[10934] = 8'b11111111;
DRAM[10935] = 8'b11111111;
DRAM[10936] = 8'b11111111;
DRAM[10937] = 8'b11111111;
DRAM[10938] = 8'b11111111;
DRAM[10939] = 8'b11111011;
DRAM[10940] = 8'b11111110;
DRAM[10941] = 8'b11111111;
DRAM[10942] = 8'b11111011;
DRAM[10943] = 8'b11101111;
DRAM[10944] = 8'b11101111;
DRAM[10945] = 8'b11110000;
DRAM[10946] = 8'b11111100;
DRAM[10947] = 8'b11110011;
DRAM[10948] = 8'b11010110;
DRAM[10949] = 8'b11001000;
DRAM[10950] = 8'b10110001;
DRAM[10951] = 8'b10001000;
DRAM[10952] = 8'b1111111;
DRAM[10953] = 8'b1111000;
DRAM[10954] = 8'b1110010;
DRAM[10955] = 8'b1110100;
DRAM[10956] = 8'b1111010;
DRAM[10957] = 8'b1111011;
DRAM[10958] = 8'b1110100;
DRAM[10959] = 8'b1101100;
DRAM[10960] = 8'b1100100;
DRAM[10961] = 8'b1100011;
DRAM[10962] = 8'b1100011;
DRAM[10963] = 8'b1100010;
DRAM[10964] = 8'b1100000;
DRAM[10965] = 8'b1011110;
DRAM[10966] = 8'b1011100;
DRAM[10967] = 8'b1011011;
DRAM[10968] = 8'b1011010;
DRAM[10969] = 8'b1011010;
DRAM[10970] = 8'b1011010;
DRAM[10971] = 8'b1011001;
DRAM[10972] = 8'b1011000;
DRAM[10973] = 8'b1010111;
DRAM[10974] = 8'b1010111;
DRAM[10975] = 8'b1010110;
DRAM[10976] = 8'b1010110;
DRAM[10977] = 8'b1010110;
DRAM[10978] = 8'b1010110;
DRAM[10979] = 8'b1010101;
DRAM[10980] = 8'b1010101;
DRAM[10981] = 8'b1010100;
DRAM[10982] = 8'b1010100;
DRAM[10983] = 8'b1010100;
DRAM[10984] = 8'b1010010;
DRAM[10985] = 8'b1010010;
DRAM[10986] = 8'b1010011;
DRAM[10987] = 8'b1010011;
DRAM[10988] = 8'b1010011;
DRAM[10989] = 8'b1010011;
DRAM[10990] = 8'b1010010;
DRAM[10991] = 8'b1010010;
DRAM[10992] = 8'b1010010;
DRAM[10993] = 8'b1010010;
DRAM[10994] = 8'b1010010;
DRAM[10995] = 8'b1010001;
DRAM[10996] = 8'b1010001;
DRAM[10997] = 8'b1010000;
DRAM[10998] = 8'b1010000;
DRAM[10999] = 8'b1010000;
DRAM[11000] = 8'b1001111;
DRAM[11001] = 8'b1001111;
DRAM[11002] = 8'b1001111;
DRAM[11003] = 8'b1001111;
DRAM[11004] = 8'b1001111;
DRAM[11005] = 8'b1001111;
DRAM[11006] = 8'b1001111;
DRAM[11007] = 8'b1001111;
DRAM[11008] = 8'b1100010;
DRAM[11009] = 8'b1100011;
DRAM[11010] = 8'b1100011;
DRAM[11011] = 8'b1100100;
DRAM[11012] = 8'b1100101;
DRAM[11013] = 8'b1100101;
DRAM[11014] = 8'b1100110;
DRAM[11015] = 8'b1100110;
DRAM[11016] = 8'b1100110;
DRAM[11017] = 8'b1100110;
DRAM[11018] = 8'b1100111;
DRAM[11019] = 8'b1101000;
DRAM[11020] = 8'b1101000;
DRAM[11021] = 8'b1101001;
DRAM[11022] = 8'b1101010;
DRAM[11023] = 8'b1101010;
DRAM[11024] = 8'b1101010;
DRAM[11025] = 8'b1101010;
DRAM[11026] = 8'b1101011;
DRAM[11027] = 8'b1101100;
DRAM[11028] = 8'b1101100;
DRAM[11029] = 8'b1101101;
DRAM[11030] = 8'b1101110;
DRAM[11031] = 8'b1101110;
DRAM[11032] = 8'b1101101;
DRAM[11033] = 8'b1101101;
DRAM[11034] = 8'b1101110;
DRAM[11035] = 8'b1101111;
DRAM[11036] = 8'b1110000;
DRAM[11037] = 8'b1110000;
DRAM[11038] = 8'b1110001;
DRAM[11039] = 8'b1110001;
DRAM[11040] = 8'b1110011;
DRAM[11041] = 8'b1110011;
DRAM[11042] = 8'b1110011;
DRAM[11043] = 8'b1110100;
DRAM[11044] = 8'b1110100;
DRAM[11045] = 8'b1110101;
DRAM[11046] = 8'b1110101;
DRAM[11047] = 8'b1110101;
DRAM[11048] = 8'b1110100;
DRAM[11049] = 8'b1110100;
DRAM[11050] = 8'b1110101;
DRAM[11051] = 8'b1110110;
DRAM[11052] = 8'b1110110;
DRAM[11053] = 8'b1110111;
DRAM[11054] = 8'b1111000;
DRAM[11055] = 8'b1111000;
DRAM[11056] = 8'b1111001;
DRAM[11057] = 8'b1111001;
DRAM[11058] = 8'b1111000;
DRAM[11059] = 8'b1111010;
DRAM[11060] = 8'b1111100;
DRAM[11061] = 8'b1111100;
DRAM[11062] = 8'b1111011;
DRAM[11063] = 8'b1111001;
DRAM[11064] = 8'b1111100;
DRAM[11065] = 8'b1111011;
DRAM[11066] = 8'b1111011;
DRAM[11067] = 8'b1111011;
DRAM[11068] = 8'b1111100;
DRAM[11069] = 8'b1111100;
DRAM[11070] = 8'b1111101;
DRAM[11071] = 8'b1111110;
DRAM[11072] = 8'b1111001;
DRAM[11073] = 8'b10000000;
DRAM[11074] = 8'b10000010;
DRAM[11075] = 8'b1111001;
DRAM[11076] = 8'b1110001;
DRAM[11077] = 8'b1110110;
DRAM[11078] = 8'b10000100;
DRAM[11079] = 8'b10010000;
DRAM[11080] = 8'b1111000;
DRAM[11081] = 8'b10001100;
DRAM[11082] = 8'b10010011;
DRAM[11083] = 8'b10010111;
DRAM[11084] = 8'b10101100;
DRAM[11085] = 8'b10111110;
DRAM[11086] = 8'b11000000;
DRAM[11087] = 8'b10111110;
DRAM[11088] = 8'b10110000;
DRAM[11089] = 8'b11001011;
DRAM[11090] = 8'b11101011;
DRAM[11091] = 8'b11111101;
DRAM[11092] = 8'b11111111;
DRAM[11093] = 8'b11111111;
DRAM[11094] = 8'b11111101;
DRAM[11095] = 8'b11111010;
DRAM[11096] = 8'b11111111;
DRAM[11097] = 8'b11111111;
DRAM[11098] = 8'b11111111;
DRAM[11099] = 8'b11111111;
DRAM[11100] = 8'b11111111;
DRAM[11101] = 8'b11111111;
DRAM[11102] = 8'b11111111;
DRAM[11103] = 8'b11111111;
DRAM[11104] = 8'b11111111;
DRAM[11105] = 8'b11111111;
DRAM[11106] = 8'b11111111;
DRAM[11107] = 8'b11111111;
DRAM[11108] = 8'b11111111;
DRAM[11109] = 8'b11111111;
DRAM[11110] = 8'b11111111;
DRAM[11111] = 8'b11111111;
DRAM[11112] = 8'b11111110;
DRAM[11113] = 8'b11111110;
DRAM[11114] = 8'b11111110;
DRAM[11115] = 8'b11111110;
DRAM[11116] = 8'b11111110;
DRAM[11117] = 8'b11111110;
DRAM[11118] = 8'b11111110;
DRAM[11119] = 8'b11111110;
DRAM[11120] = 8'b11111110;
DRAM[11121] = 8'b11111110;
DRAM[11122] = 8'b11111110;
DRAM[11123] = 8'b11111110;
DRAM[11124] = 8'b11111110;
DRAM[11125] = 8'b11111110;
DRAM[11126] = 8'b11111110;
DRAM[11127] = 8'b11111110;
DRAM[11128] = 8'b11111110;
DRAM[11129] = 8'b11111110;
DRAM[11130] = 8'b11111110;
DRAM[11131] = 8'b11111111;
DRAM[11132] = 8'b11111111;
DRAM[11133] = 8'b11111111;
DRAM[11134] = 8'b11111111;
DRAM[11135] = 8'b11111111;
DRAM[11136] = 8'b11111111;
DRAM[11137] = 8'b11111111;
DRAM[11138] = 8'b11111111;
DRAM[11139] = 8'b11111111;
DRAM[11140] = 8'b11111111;
DRAM[11141] = 8'b11111111;
DRAM[11142] = 8'b11111111;
DRAM[11143] = 8'b11111111;
DRAM[11144] = 8'b11111111;
DRAM[11145] = 8'b11111111;
DRAM[11146] = 8'b11111111;
DRAM[11147] = 8'b11111111;
DRAM[11148] = 8'b11111111;
DRAM[11149] = 8'b11111111;
DRAM[11150] = 8'b11111111;
DRAM[11151] = 8'b11111111;
DRAM[11152] = 8'b11111110;
DRAM[11153] = 8'b11111110;
DRAM[11154] = 8'b11111110;
DRAM[11155] = 8'b11111110;
DRAM[11156] = 8'b11111110;
DRAM[11157] = 8'b11111110;
DRAM[11158] = 8'b11111110;
DRAM[11159] = 8'b11111110;
DRAM[11160] = 8'b11111110;
DRAM[11161] = 8'b11111110;
DRAM[11162] = 8'b11111110;
DRAM[11163] = 8'b11111111;
DRAM[11164] = 8'b11111111;
DRAM[11165] = 8'b11111111;
DRAM[11166] = 8'b11111111;
DRAM[11167] = 8'b11111111;
DRAM[11168] = 8'b11111110;
DRAM[11169] = 8'b11111110;
DRAM[11170] = 8'b11111110;
DRAM[11171] = 8'b11111110;
DRAM[11172] = 8'b11111110;
DRAM[11173] = 8'b11111110;
DRAM[11174] = 8'b11111110;
DRAM[11175] = 8'b11111110;
DRAM[11176] = 8'b11111101;
DRAM[11177] = 8'b11111101;
DRAM[11178] = 8'b11111101;
DRAM[11179] = 8'b11111110;
DRAM[11180] = 8'b11111110;
DRAM[11181] = 8'b11111111;
DRAM[11182] = 8'b11111111;
DRAM[11183] = 8'b11111111;
DRAM[11184] = 8'b11111111;
DRAM[11185] = 8'b11111111;
DRAM[11186] = 8'b11111111;
DRAM[11187] = 8'b11111111;
DRAM[11188] = 8'b11111111;
DRAM[11189] = 8'b11111111;
DRAM[11190] = 8'b11111111;
DRAM[11191] = 8'b11111111;
DRAM[11192] = 8'b11111111;
DRAM[11193] = 8'b11111111;
DRAM[11194] = 8'b11111110;
DRAM[11195] = 8'b11111011;
DRAM[11196] = 8'b11111111;
DRAM[11197] = 8'b11111111;
DRAM[11198] = 8'b11111111;
DRAM[11199] = 8'b11111000;
DRAM[11200] = 8'b11111111;
DRAM[11201] = 8'b11111101;
DRAM[11202] = 8'b11111111;
DRAM[11203] = 8'b11111111;
DRAM[11204] = 8'b11111001;
DRAM[11205] = 8'b11110110;
DRAM[11206] = 8'b11011001;
DRAM[11207] = 8'b10101001;
DRAM[11208] = 8'b10101101;
DRAM[11209] = 8'b10100101;
DRAM[11210] = 8'b10011001;
DRAM[11211] = 8'b10001110;
DRAM[11212] = 8'b10000011;
DRAM[11213] = 8'b1111001;
DRAM[11214] = 8'b1101110;
DRAM[11215] = 8'b1100110;
DRAM[11216] = 8'b1100101;
DRAM[11217] = 8'b1100101;
DRAM[11218] = 8'b1100100;
DRAM[11219] = 8'b1100011;
DRAM[11220] = 8'b1100011;
DRAM[11221] = 8'b1100001;
DRAM[11222] = 8'b1011110;
DRAM[11223] = 8'b1011100;
DRAM[11224] = 8'b1011011;
DRAM[11225] = 8'b1011011;
DRAM[11226] = 8'b1011010;
DRAM[11227] = 8'b1011001;
DRAM[11228] = 8'b1011000;
DRAM[11229] = 8'b1011000;
DRAM[11230] = 8'b1010111;
DRAM[11231] = 8'b1010111;
DRAM[11232] = 8'b1010110;
DRAM[11233] = 8'b1010110;
DRAM[11234] = 8'b1010110;
DRAM[11235] = 8'b1010101;
DRAM[11236] = 8'b1010101;
DRAM[11237] = 8'b1010100;
DRAM[11238] = 8'b1010100;
DRAM[11239] = 8'b1010100;
DRAM[11240] = 8'b1010010;
DRAM[11241] = 8'b1010010;
DRAM[11242] = 8'b1010011;
DRAM[11243] = 8'b1010100;
DRAM[11244] = 8'b1010100;
DRAM[11245] = 8'b1010011;
DRAM[11246] = 8'b1010010;
DRAM[11247] = 8'b1010010;
DRAM[11248] = 8'b1010010;
DRAM[11249] = 8'b1010010;
DRAM[11250] = 8'b1010010;
DRAM[11251] = 8'b1010001;
DRAM[11252] = 8'b1010001;
DRAM[11253] = 8'b1010000;
DRAM[11254] = 8'b1010000;
DRAM[11255] = 8'b1010000;
DRAM[11256] = 8'b1001110;
DRAM[11257] = 8'b1001110;
DRAM[11258] = 8'b1001110;
DRAM[11259] = 8'b1001110;
DRAM[11260] = 8'b1001110;
DRAM[11261] = 8'b1001110;
DRAM[11262] = 8'b1001110;
DRAM[11263] = 8'b1001110;
DRAM[11264] = 8'b1100100;
DRAM[11265] = 8'b1100100;
DRAM[11266] = 8'b1100101;
DRAM[11267] = 8'b1100101;
DRAM[11268] = 8'b1100110;
DRAM[11269] = 8'b1100111;
DRAM[11270] = 8'b1100111;
DRAM[11271] = 8'b1101000;
DRAM[11272] = 8'b1100110;
DRAM[11273] = 8'b1100110;
DRAM[11274] = 8'b1100111;
DRAM[11275] = 8'b1101000;
DRAM[11276] = 8'b1101000;
DRAM[11277] = 8'b1101001;
DRAM[11278] = 8'b1101010;
DRAM[11279] = 8'b1101010;
DRAM[11280] = 8'b1101010;
DRAM[11281] = 8'b1101010;
DRAM[11282] = 8'b1101011;
DRAM[11283] = 8'b1101100;
DRAM[11284] = 8'b1101100;
DRAM[11285] = 8'b1101101;
DRAM[11286] = 8'b1101110;
DRAM[11287] = 8'b1101110;
DRAM[11288] = 8'b1101101;
DRAM[11289] = 8'b1101101;
DRAM[11290] = 8'b1101110;
DRAM[11291] = 8'b1101110;
DRAM[11292] = 8'b1101111;
DRAM[11293] = 8'b1110000;
DRAM[11294] = 8'b1110001;
DRAM[11295] = 8'b1110001;
DRAM[11296] = 8'b1110011;
DRAM[11297] = 8'b1110011;
DRAM[11298] = 8'b1110011;
DRAM[11299] = 8'b1110100;
DRAM[11300] = 8'b1110100;
DRAM[11301] = 8'b1110101;
DRAM[11302] = 8'b1110101;
DRAM[11303] = 8'b1110101;
DRAM[11304] = 8'b1110100;
DRAM[11305] = 8'b1110100;
DRAM[11306] = 8'b1110101;
DRAM[11307] = 8'b1110110;
DRAM[11308] = 8'b1110110;
DRAM[11309] = 8'b1110111;
DRAM[11310] = 8'b1111000;
DRAM[11311] = 8'b1111000;
DRAM[11312] = 8'b1111001;
DRAM[11313] = 8'b1111001;
DRAM[11314] = 8'b1111000;
DRAM[11315] = 8'b1111010;
DRAM[11316] = 8'b1111100;
DRAM[11317] = 8'b1111100;
DRAM[11318] = 8'b1111011;
DRAM[11319] = 8'b1111001;
DRAM[11320] = 8'b1111010;
DRAM[11321] = 8'b1111010;
DRAM[11322] = 8'b1111011;
DRAM[11323] = 8'b1111100;
DRAM[11324] = 8'b1111110;
DRAM[11325] = 8'b10000000;
DRAM[11326] = 8'b10000010;
DRAM[11327] = 8'b10000100;
DRAM[11328] = 8'b1111100;
DRAM[11329] = 8'b10000100;
DRAM[11330] = 8'b10001001;
DRAM[11331] = 8'b10000111;
DRAM[11332] = 8'b10001010;
DRAM[11333] = 8'b10010101;
DRAM[11334] = 8'b10100001;
DRAM[11335] = 8'b10100111;
DRAM[11336] = 8'b10100100;
DRAM[11337] = 8'b10011111;
DRAM[11338] = 8'b10100100;
DRAM[11339] = 8'b10111111;
DRAM[11340] = 8'b11010101;
DRAM[11341] = 8'b11010001;
DRAM[11342] = 8'b11010110;
DRAM[11343] = 8'b11101111;
DRAM[11344] = 8'b11110100;
DRAM[11345] = 8'b11110111;
DRAM[11346] = 8'b11110111;
DRAM[11347] = 8'b11110100;
DRAM[11348] = 8'b11110101;
DRAM[11349] = 8'b11111010;
DRAM[11350] = 8'b11111111;
DRAM[11351] = 8'b11111111;
DRAM[11352] = 8'b11111111;
DRAM[11353] = 8'b11111111;
DRAM[11354] = 8'b11111111;
DRAM[11355] = 8'b11111111;
DRAM[11356] = 8'b11111111;
DRAM[11357] = 8'b11111111;
DRAM[11358] = 8'b11111111;
DRAM[11359] = 8'b11111111;
DRAM[11360] = 8'b11111111;
DRAM[11361] = 8'b11111111;
DRAM[11362] = 8'b11111111;
DRAM[11363] = 8'b11111111;
DRAM[11364] = 8'b11111111;
DRAM[11365] = 8'b11111111;
DRAM[11366] = 8'b11111111;
DRAM[11367] = 8'b11111111;
DRAM[11368] = 8'b11111110;
DRAM[11369] = 8'b11111110;
DRAM[11370] = 8'b11111110;
DRAM[11371] = 8'b11111110;
DRAM[11372] = 8'b11111110;
DRAM[11373] = 8'b11111110;
DRAM[11374] = 8'b11111110;
DRAM[11375] = 8'b11111110;
DRAM[11376] = 8'b11111110;
DRAM[11377] = 8'b11111110;
DRAM[11378] = 8'b11111110;
DRAM[11379] = 8'b11111110;
DRAM[11380] = 8'b11111110;
DRAM[11381] = 8'b11111110;
DRAM[11382] = 8'b11111110;
DRAM[11383] = 8'b11111110;
DRAM[11384] = 8'b11111110;
DRAM[11385] = 8'b11111110;
DRAM[11386] = 8'b11111110;
DRAM[11387] = 8'b11111111;
DRAM[11388] = 8'b11111111;
DRAM[11389] = 8'b11111111;
DRAM[11390] = 8'b11111111;
DRAM[11391] = 8'b11111111;
DRAM[11392] = 8'b11111111;
DRAM[11393] = 8'b11111111;
DRAM[11394] = 8'b11111111;
DRAM[11395] = 8'b11111111;
DRAM[11396] = 8'b11111111;
DRAM[11397] = 8'b11111111;
DRAM[11398] = 8'b11111111;
DRAM[11399] = 8'b11111111;
DRAM[11400] = 8'b11111111;
DRAM[11401] = 8'b11111111;
DRAM[11402] = 8'b11111111;
DRAM[11403] = 8'b11111111;
DRAM[11404] = 8'b11111111;
DRAM[11405] = 8'b11111111;
DRAM[11406] = 8'b11111111;
DRAM[11407] = 8'b11111111;
DRAM[11408] = 8'b11111110;
DRAM[11409] = 8'b11111110;
DRAM[11410] = 8'b11111110;
DRAM[11411] = 8'b11111110;
DRAM[11412] = 8'b11111110;
DRAM[11413] = 8'b11111110;
DRAM[11414] = 8'b11111110;
DRAM[11415] = 8'b11111110;
DRAM[11416] = 8'b11111110;
DRAM[11417] = 8'b11111110;
DRAM[11418] = 8'b11111110;
DRAM[11419] = 8'b11111111;
DRAM[11420] = 8'b11111111;
DRAM[11421] = 8'b11111111;
DRAM[11422] = 8'b11111111;
DRAM[11423] = 8'b11111111;
DRAM[11424] = 8'b11111110;
DRAM[11425] = 8'b11111110;
DRAM[11426] = 8'b11111110;
DRAM[11427] = 8'b11111110;
DRAM[11428] = 8'b11111110;
DRAM[11429] = 8'b11111110;
DRAM[11430] = 8'b11111110;
DRAM[11431] = 8'b11111110;
DRAM[11432] = 8'b11111101;
DRAM[11433] = 8'b11111101;
DRAM[11434] = 8'b11111101;
DRAM[11435] = 8'b11111110;
DRAM[11436] = 8'b11111110;
DRAM[11437] = 8'b11111111;
DRAM[11438] = 8'b11111111;
DRAM[11439] = 8'b11111111;
DRAM[11440] = 8'b11111111;
DRAM[11441] = 8'b11111111;
DRAM[11442] = 8'b11111111;
DRAM[11443] = 8'b11111111;
DRAM[11444] = 8'b11111111;
DRAM[11445] = 8'b11111111;
DRAM[11446] = 8'b11111111;
DRAM[11447] = 8'b11111111;
DRAM[11448] = 8'b11111111;
DRAM[11449] = 8'b11111110;
DRAM[11450] = 8'b11111100;
DRAM[11451] = 8'b11111011;
DRAM[11452] = 8'b11111110;
DRAM[11453] = 8'b11111111;
DRAM[11454] = 8'b11111111;
DRAM[11455] = 8'b11111101;
DRAM[11456] = 8'b11111010;
DRAM[11457] = 8'b11111010;
DRAM[11458] = 8'b11111101;
DRAM[11459] = 8'b11111011;
DRAM[11460] = 8'b11110101;
DRAM[11461] = 8'b11111000;
DRAM[11462] = 8'b11111011;
DRAM[11463] = 8'b11110111;
DRAM[11464] = 8'b11100110;
DRAM[11465] = 8'b11011001;
DRAM[11466] = 8'b11000001;
DRAM[11467] = 8'b10100011;
DRAM[11468] = 8'b10001000;
DRAM[11469] = 8'b1110110;
DRAM[11470] = 8'b1101111;
DRAM[11471] = 8'b1101110;
DRAM[11472] = 8'b1101000;
DRAM[11473] = 8'b1100101;
DRAM[11474] = 8'b1100011;
DRAM[11475] = 8'b1100011;
DRAM[11476] = 8'b1100011;
DRAM[11477] = 8'b1100010;
DRAM[11478] = 8'b1011111;
DRAM[11479] = 8'b1011100;
DRAM[11480] = 8'b1011011;
DRAM[11481] = 8'b1011011;
DRAM[11482] = 8'b1011010;
DRAM[11483] = 8'b1011010;
DRAM[11484] = 8'b1011001;
DRAM[11485] = 8'b1011000;
DRAM[11486] = 8'b1010111;
DRAM[11487] = 8'b1010111;
DRAM[11488] = 8'b1010110;
DRAM[11489] = 8'b1010110;
DRAM[11490] = 8'b1010110;
DRAM[11491] = 8'b1010101;
DRAM[11492] = 8'b1010101;
DRAM[11493] = 8'b1010100;
DRAM[11494] = 8'b1010100;
DRAM[11495] = 8'b1010100;
DRAM[11496] = 8'b1010010;
DRAM[11497] = 8'b1010011;
DRAM[11498] = 8'b1010100;
DRAM[11499] = 8'b1010100;
DRAM[11500] = 8'b1010100;
DRAM[11501] = 8'b1010100;
DRAM[11502] = 8'b1010011;
DRAM[11503] = 8'b1010010;
DRAM[11504] = 8'b1010010;
DRAM[11505] = 8'b1010010;
DRAM[11506] = 8'b1010010;
DRAM[11507] = 8'b1010001;
DRAM[11508] = 8'b1010001;
DRAM[11509] = 8'b1010000;
DRAM[11510] = 8'b1010000;
DRAM[11511] = 8'b1010000;
DRAM[11512] = 8'b1001110;
DRAM[11513] = 8'b1001110;
DRAM[11514] = 8'b1001110;
DRAM[11515] = 8'b1001110;
DRAM[11516] = 8'b1001110;
DRAM[11517] = 8'b1001110;
DRAM[11518] = 8'b1001110;
DRAM[11519] = 8'b1001110;
DRAM[11520] = 8'b1100100;
DRAM[11521] = 8'b1100100;
DRAM[11522] = 8'b1100101;
DRAM[11523] = 8'b1100110;
DRAM[11524] = 8'b1100111;
DRAM[11525] = 8'b1100111;
DRAM[11526] = 8'b1101000;
DRAM[11527] = 8'b1101000;
DRAM[11528] = 8'b1100110;
DRAM[11529] = 8'b1100110;
DRAM[11530] = 8'b1100111;
DRAM[11531] = 8'b1101000;
DRAM[11532] = 8'b1101000;
DRAM[11533] = 8'b1101001;
DRAM[11534] = 8'b1101010;
DRAM[11535] = 8'b1101010;
DRAM[11536] = 8'b1101010;
DRAM[11537] = 8'b1101010;
DRAM[11538] = 8'b1101011;
DRAM[11539] = 8'b1101100;
DRAM[11540] = 8'b1101100;
DRAM[11541] = 8'b1101101;
DRAM[11542] = 8'b1101110;
DRAM[11543] = 8'b1101110;
DRAM[11544] = 8'b1101110;
DRAM[11545] = 8'b1101110;
DRAM[11546] = 8'b1101101;
DRAM[11547] = 8'b1101110;
DRAM[11548] = 8'b1101111;
DRAM[11549] = 8'b1110000;
DRAM[11550] = 8'b1110001;
DRAM[11551] = 8'b1110010;
DRAM[11552] = 8'b1110011;
DRAM[11553] = 8'b1110011;
DRAM[11554] = 8'b1110011;
DRAM[11555] = 8'b1110100;
DRAM[11556] = 8'b1110100;
DRAM[11557] = 8'b1110101;
DRAM[11558] = 8'b1110101;
DRAM[11559] = 8'b1110101;
DRAM[11560] = 8'b1110100;
DRAM[11561] = 8'b1110100;
DRAM[11562] = 8'b1110101;
DRAM[11563] = 8'b1110110;
DRAM[11564] = 8'b1110110;
DRAM[11565] = 8'b1110111;
DRAM[11566] = 8'b1111000;
DRAM[11567] = 8'b1111000;
DRAM[11568] = 8'b1111001;
DRAM[11569] = 8'b1111001;
DRAM[11570] = 8'b1111000;
DRAM[11571] = 8'b1111010;
DRAM[11572] = 8'b1111100;
DRAM[11573] = 8'b1111100;
DRAM[11574] = 8'b1111011;
DRAM[11575] = 8'b1111001;
DRAM[11576] = 8'b1111001;
DRAM[11577] = 8'b1111001;
DRAM[11578] = 8'b1111010;
DRAM[11579] = 8'b1111101;
DRAM[11580] = 8'b10000001;
DRAM[11581] = 8'b10000101;
DRAM[11582] = 8'b10001001;
DRAM[11583] = 8'b10001100;
DRAM[11584] = 8'b1111011;
DRAM[11585] = 8'b1111101;
DRAM[11586] = 8'b10000001;
DRAM[11587] = 8'b10001110;
DRAM[11588] = 8'b10101011;
DRAM[11589] = 8'b11001010;
DRAM[11590] = 8'b11010111;
DRAM[11591] = 8'b11010110;
DRAM[11592] = 8'b11111001;
DRAM[11593] = 8'b11110111;
DRAM[11594] = 8'b11110001;
DRAM[11595] = 8'b11110110;
DRAM[11596] = 8'b11111111;
DRAM[11597] = 8'b11111010;
DRAM[11598] = 8'b11110111;
DRAM[11599] = 8'b11111111;
DRAM[11600] = 8'b11111011;
DRAM[11601] = 8'b11111101;
DRAM[11602] = 8'b11111101;
DRAM[11603] = 8'b11111100;
DRAM[11604] = 8'b11111110;
DRAM[11605] = 8'b11111111;
DRAM[11606] = 8'b11111100;
DRAM[11607] = 8'b11110110;
DRAM[11608] = 8'b11111110;
DRAM[11609] = 8'b11111110;
DRAM[11610] = 8'b11111101;
DRAM[11611] = 8'b11111110;
DRAM[11612] = 8'b11111111;
DRAM[11613] = 8'b11111111;
DRAM[11614] = 8'b11111111;
DRAM[11615] = 8'b11111111;
DRAM[11616] = 8'b11111111;
DRAM[11617] = 8'b11111111;
DRAM[11618] = 8'b11111111;
DRAM[11619] = 8'b11111111;
DRAM[11620] = 8'b11111111;
DRAM[11621] = 8'b11111111;
DRAM[11622] = 8'b11111111;
DRAM[11623] = 8'b11111111;
DRAM[11624] = 8'b11111110;
DRAM[11625] = 8'b11111110;
DRAM[11626] = 8'b11111110;
DRAM[11627] = 8'b11111110;
DRAM[11628] = 8'b11111110;
DRAM[11629] = 8'b11111110;
DRAM[11630] = 8'b11111110;
DRAM[11631] = 8'b11111110;
DRAM[11632] = 8'b11111110;
DRAM[11633] = 8'b11111110;
DRAM[11634] = 8'b11111110;
DRAM[11635] = 8'b11111110;
DRAM[11636] = 8'b11111110;
DRAM[11637] = 8'b11111110;
DRAM[11638] = 8'b11111110;
DRAM[11639] = 8'b11111110;
DRAM[11640] = 8'b11111110;
DRAM[11641] = 8'b11111110;
DRAM[11642] = 8'b11111110;
DRAM[11643] = 8'b11111111;
DRAM[11644] = 8'b11111111;
DRAM[11645] = 8'b11111111;
DRAM[11646] = 8'b11111111;
DRAM[11647] = 8'b11111111;
DRAM[11648] = 8'b11111111;
DRAM[11649] = 8'b11111111;
DRAM[11650] = 8'b11111111;
DRAM[11651] = 8'b11111111;
DRAM[11652] = 8'b11111111;
DRAM[11653] = 8'b11111111;
DRAM[11654] = 8'b11111111;
DRAM[11655] = 8'b11111111;
DRAM[11656] = 8'b11111111;
DRAM[11657] = 8'b11111111;
DRAM[11658] = 8'b11111111;
DRAM[11659] = 8'b11111111;
DRAM[11660] = 8'b11111111;
DRAM[11661] = 8'b11111111;
DRAM[11662] = 8'b11111111;
DRAM[11663] = 8'b11111111;
DRAM[11664] = 8'b11111111;
DRAM[11665] = 8'b11111111;
DRAM[11666] = 8'b11111110;
DRAM[11667] = 8'b11111110;
DRAM[11668] = 8'b11111110;
DRAM[11669] = 8'b11111110;
DRAM[11670] = 8'b11111101;
DRAM[11671] = 8'b11111101;
DRAM[11672] = 8'b11111110;
DRAM[11673] = 8'b11111110;
DRAM[11674] = 8'b11111110;
DRAM[11675] = 8'b11111111;
DRAM[11676] = 8'b11111111;
DRAM[11677] = 8'b11111111;
DRAM[11678] = 8'b11111111;
DRAM[11679] = 8'b11111111;
DRAM[11680] = 8'b11111110;
DRAM[11681] = 8'b11111110;
DRAM[11682] = 8'b11111110;
DRAM[11683] = 8'b11111110;
DRAM[11684] = 8'b11111110;
DRAM[11685] = 8'b11111110;
DRAM[11686] = 8'b11111110;
DRAM[11687] = 8'b11111110;
DRAM[11688] = 8'b11111101;
DRAM[11689] = 8'b11111101;
DRAM[11690] = 8'b11111101;
DRAM[11691] = 8'b11111110;
DRAM[11692] = 8'b11111110;
DRAM[11693] = 8'b11111111;
DRAM[11694] = 8'b11111111;
DRAM[11695] = 8'b11111111;
DRAM[11696] = 8'b11111111;
DRAM[11697] = 8'b11111111;
DRAM[11698] = 8'b11111111;
DRAM[11699] = 8'b11111111;
DRAM[11700] = 8'b11111111;
DRAM[11701] = 8'b11111111;
DRAM[11702] = 8'b11111111;
DRAM[11703] = 8'b11111111;
DRAM[11704] = 8'b11111111;
DRAM[11705] = 8'b11111101;
DRAM[11706] = 8'b11111100;
DRAM[11707] = 8'b11111011;
DRAM[11708] = 8'b11111101;
DRAM[11709] = 8'b11111111;
DRAM[11710] = 8'b11111111;
DRAM[11711] = 8'b11111110;
DRAM[11712] = 8'b11111111;
DRAM[11713] = 8'b11111100;
DRAM[11714] = 8'b11111010;
DRAM[11715] = 8'b11111100;
DRAM[11716] = 8'b11111101;
DRAM[11717] = 8'b11111011;
DRAM[11718] = 8'b11111110;
DRAM[11719] = 8'b11111111;
DRAM[11720] = 8'b11110001;
DRAM[11721] = 8'b11100100;
DRAM[11722] = 8'b11001100;
DRAM[11723] = 8'b10101101;
DRAM[11724] = 8'b10010011;
DRAM[11725] = 8'b10000110;
DRAM[11726] = 8'b10000100;
DRAM[11727] = 8'b10000111;
DRAM[11728] = 8'b1101010;
DRAM[11729] = 8'b1100110;
DRAM[11730] = 8'b1100010;
DRAM[11731] = 8'b1100001;
DRAM[11732] = 8'b1100010;
DRAM[11733] = 8'b1100011;
DRAM[11734] = 8'b1100000;
DRAM[11735] = 8'b1011101;
DRAM[11736] = 8'b1011100;
DRAM[11737] = 8'b1011011;
DRAM[11738] = 8'b1011011;
DRAM[11739] = 8'b1011010;
DRAM[11740] = 8'b1011001;
DRAM[11741] = 8'b1011000;
DRAM[11742] = 8'b1011000;
DRAM[11743] = 8'b1011000;
DRAM[11744] = 8'b1010110;
DRAM[11745] = 8'b1010110;
DRAM[11746] = 8'b1010110;
DRAM[11747] = 8'b1010101;
DRAM[11748] = 8'b1010101;
DRAM[11749] = 8'b1010100;
DRAM[11750] = 8'b1010100;
DRAM[11751] = 8'b1010100;
DRAM[11752] = 8'b1010011;
DRAM[11753] = 8'b1010011;
DRAM[11754] = 8'b1010100;
DRAM[11755] = 8'b1010100;
DRAM[11756] = 8'b1010100;
DRAM[11757] = 8'b1010100;
DRAM[11758] = 8'b1010011;
DRAM[11759] = 8'b1010011;
DRAM[11760] = 8'b1010010;
DRAM[11761] = 8'b1010010;
DRAM[11762] = 8'b1010010;
DRAM[11763] = 8'b1010001;
DRAM[11764] = 8'b1010001;
DRAM[11765] = 8'b1010000;
DRAM[11766] = 8'b1010000;
DRAM[11767] = 8'b1010000;
DRAM[11768] = 8'b1001111;
DRAM[11769] = 8'b1001111;
DRAM[11770] = 8'b1001111;
DRAM[11771] = 8'b1001111;
DRAM[11772] = 8'b1001111;
DRAM[11773] = 8'b1001111;
DRAM[11774] = 8'b1001111;
DRAM[11775] = 8'b1001111;
DRAM[11776] = 8'b1100011;
DRAM[11777] = 8'b1100011;
DRAM[11778] = 8'b1100100;
DRAM[11779] = 8'b1100101;
DRAM[11780] = 8'b1100110;
DRAM[11781] = 8'b1100110;
DRAM[11782] = 8'b1100111;
DRAM[11783] = 8'b1100111;
DRAM[11784] = 8'b1100110;
DRAM[11785] = 8'b1100110;
DRAM[11786] = 8'b1100111;
DRAM[11787] = 8'b1101000;
DRAM[11788] = 8'b1101000;
DRAM[11789] = 8'b1101001;
DRAM[11790] = 8'b1101010;
DRAM[11791] = 8'b1101010;
DRAM[11792] = 8'b1101010;
DRAM[11793] = 8'b1101010;
DRAM[11794] = 8'b1101011;
DRAM[11795] = 8'b1101100;
DRAM[11796] = 8'b1101100;
DRAM[11797] = 8'b1101101;
DRAM[11798] = 8'b1101110;
DRAM[11799] = 8'b1101110;
DRAM[11800] = 8'b1101110;
DRAM[11801] = 8'b1101110;
DRAM[11802] = 8'b1101101;
DRAM[11803] = 8'b1101101;
DRAM[11804] = 8'b1101110;
DRAM[11805] = 8'b1110000;
DRAM[11806] = 8'b1110001;
DRAM[11807] = 8'b1110010;
DRAM[11808] = 8'b1110011;
DRAM[11809] = 8'b1110011;
DRAM[11810] = 8'b1110011;
DRAM[11811] = 8'b1110100;
DRAM[11812] = 8'b1110100;
DRAM[11813] = 8'b1110101;
DRAM[11814] = 8'b1110101;
DRAM[11815] = 8'b1110101;
DRAM[11816] = 8'b1110100;
DRAM[11817] = 8'b1110100;
DRAM[11818] = 8'b1110101;
DRAM[11819] = 8'b1110110;
DRAM[11820] = 8'b1110110;
DRAM[11821] = 8'b1110111;
DRAM[11822] = 8'b1111000;
DRAM[11823] = 8'b1111000;
DRAM[11824] = 8'b1111001;
DRAM[11825] = 8'b1111001;
DRAM[11826] = 8'b1111000;
DRAM[11827] = 8'b1111010;
DRAM[11828] = 8'b1111100;
DRAM[11829] = 8'b1111100;
DRAM[11830] = 8'b1111011;
DRAM[11831] = 8'b1111001;
DRAM[11832] = 8'b1111010;
DRAM[11833] = 8'b1111010;
DRAM[11834] = 8'b1111010;
DRAM[11835] = 8'b1111011;
DRAM[11836] = 8'b1111110;
DRAM[11837] = 8'b10000010;
DRAM[11838] = 8'b10000110;
DRAM[11839] = 8'b10001000;
DRAM[11840] = 8'b10010010;
DRAM[11841] = 8'b10001110;
DRAM[11842] = 8'b10000110;
DRAM[11843] = 8'b10001000;
DRAM[11844] = 8'b10100101;
DRAM[11845] = 8'b11010011;
DRAM[11846] = 8'b11110110;
DRAM[11847] = 8'b11111111;
DRAM[11848] = 8'b11101010;
DRAM[11849] = 8'b11111001;
DRAM[11850] = 8'b11110100;
DRAM[11851] = 8'b11101000;
DRAM[11852] = 8'b11110001;
DRAM[11853] = 8'b11111101;
DRAM[11854] = 8'b11111010;
DRAM[11855] = 8'b11110100;
DRAM[11856] = 8'b11111010;
DRAM[11857] = 8'b11111001;
DRAM[11858] = 8'b11110101;
DRAM[11859] = 8'b11110001;
DRAM[11860] = 8'b11110011;
DRAM[11861] = 8'b11111100;
DRAM[11862] = 8'b11111111;
DRAM[11863] = 8'b11111111;
DRAM[11864] = 8'b11111110;
DRAM[11865] = 8'b11111110;
DRAM[11866] = 8'b11111110;
DRAM[11867] = 8'b11111111;
DRAM[11868] = 8'b11111111;
DRAM[11869] = 8'b11111111;
DRAM[11870] = 8'b11111111;
DRAM[11871] = 8'b11111111;
DRAM[11872] = 8'b11111111;
DRAM[11873] = 8'b11111111;
DRAM[11874] = 8'b11111111;
DRAM[11875] = 8'b11111111;
DRAM[11876] = 8'b11111111;
DRAM[11877] = 8'b11111111;
DRAM[11878] = 8'b11111111;
DRAM[11879] = 8'b11111111;
DRAM[11880] = 8'b11111110;
DRAM[11881] = 8'b11111110;
DRAM[11882] = 8'b11111110;
DRAM[11883] = 8'b11111110;
DRAM[11884] = 8'b11111110;
DRAM[11885] = 8'b11111110;
DRAM[11886] = 8'b11111110;
DRAM[11887] = 8'b11111110;
DRAM[11888] = 8'b11111110;
DRAM[11889] = 8'b11111110;
DRAM[11890] = 8'b11111110;
DRAM[11891] = 8'b11111110;
DRAM[11892] = 8'b11111110;
DRAM[11893] = 8'b11111110;
DRAM[11894] = 8'b11111110;
DRAM[11895] = 8'b11111110;
DRAM[11896] = 8'b11111110;
DRAM[11897] = 8'b11111110;
DRAM[11898] = 8'b11111110;
DRAM[11899] = 8'b11111111;
DRAM[11900] = 8'b11111111;
DRAM[11901] = 8'b11111111;
DRAM[11902] = 8'b11111111;
DRAM[11903] = 8'b11111111;
DRAM[11904] = 8'b11111111;
DRAM[11905] = 8'b11111111;
DRAM[11906] = 8'b11111111;
DRAM[11907] = 8'b11111111;
DRAM[11908] = 8'b11111111;
DRAM[11909] = 8'b11111111;
DRAM[11910] = 8'b11111111;
DRAM[11911] = 8'b11111111;
DRAM[11912] = 8'b11111111;
DRAM[11913] = 8'b11111111;
DRAM[11914] = 8'b11111111;
DRAM[11915] = 8'b11111111;
DRAM[11916] = 8'b11111111;
DRAM[11917] = 8'b11111111;
DRAM[11918] = 8'b11111111;
DRAM[11919] = 8'b11111111;
DRAM[11920] = 8'b11111111;
DRAM[11921] = 8'b11111111;
DRAM[11922] = 8'b11111111;
DRAM[11923] = 8'b11111110;
DRAM[11924] = 8'b11111110;
DRAM[11925] = 8'b11111101;
DRAM[11926] = 8'b11111101;
DRAM[11927] = 8'b11111101;
DRAM[11928] = 8'b11111110;
DRAM[11929] = 8'b11111110;
DRAM[11930] = 8'b11111110;
DRAM[11931] = 8'b11111111;
DRAM[11932] = 8'b11111111;
DRAM[11933] = 8'b11111111;
DRAM[11934] = 8'b11111111;
DRAM[11935] = 8'b11111111;
DRAM[11936] = 8'b11111110;
DRAM[11937] = 8'b11111110;
DRAM[11938] = 8'b11111110;
DRAM[11939] = 8'b11111110;
DRAM[11940] = 8'b11111110;
DRAM[11941] = 8'b11111110;
DRAM[11942] = 8'b11111110;
DRAM[11943] = 8'b11111110;
DRAM[11944] = 8'b11111101;
DRAM[11945] = 8'b11111101;
DRAM[11946] = 8'b11111101;
DRAM[11947] = 8'b11111110;
DRAM[11948] = 8'b11111110;
DRAM[11949] = 8'b11111111;
DRAM[11950] = 8'b11111111;
DRAM[11951] = 8'b11111111;
DRAM[11952] = 8'b11111111;
DRAM[11953] = 8'b11111111;
DRAM[11954] = 8'b11111111;
DRAM[11955] = 8'b11111111;
DRAM[11956] = 8'b11111111;
DRAM[11957] = 8'b11111111;
DRAM[11958] = 8'b11111111;
DRAM[11959] = 8'b11111111;
DRAM[11960] = 8'b11111111;
DRAM[11961] = 8'b11111110;
DRAM[11962] = 8'b11111101;
DRAM[11963] = 8'b11111101;
DRAM[11964] = 8'b11111110;
DRAM[11965] = 8'b11111101;
DRAM[11966] = 8'b11111101;
DRAM[11967] = 8'b11111101;
DRAM[11968] = 8'b11111111;
DRAM[11969] = 8'b11111111;
DRAM[11970] = 8'b11111010;
DRAM[11971] = 8'b11111110;
DRAM[11972] = 8'b11111111;
DRAM[11973] = 8'b11111111;
DRAM[11974] = 8'b11110110;
DRAM[11975] = 8'b11110000;
DRAM[11976] = 8'b11111101;
DRAM[11977] = 8'b11110100;
DRAM[11978] = 8'b11100100;
DRAM[11979] = 8'b11010000;
DRAM[11980] = 8'b10111001;
DRAM[11981] = 8'b10100001;
DRAM[11982] = 8'b10001101;
DRAM[11983] = 8'b10000001;
DRAM[11984] = 8'b1101100;
DRAM[11985] = 8'b1100110;
DRAM[11986] = 8'b1100000;
DRAM[11987] = 8'b1011110;
DRAM[11988] = 8'b1100001;
DRAM[11989] = 8'b1100010;
DRAM[11990] = 8'b1100001;
DRAM[11991] = 8'b1011110;
DRAM[11992] = 8'b1011100;
DRAM[11993] = 8'b1011100;
DRAM[11994] = 8'b1011011;
DRAM[11995] = 8'b1011010;
DRAM[11996] = 8'b1011001;
DRAM[11997] = 8'b1011001;
DRAM[11998] = 8'b1011000;
DRAM[11999] = 8'b1011000;
DRAM[12000] = 8'b1010110;
DRAM[12001] = 8'b1010110;
DRAM[12002] = 8'b1010110;
DRAM[12003] = 8'b1010101;
DRAM[12004] = 8'b1010101;
DRAM[12005] = 8'b1010100;
DRAM[12006] = 8'b1010100;
DRAM[12007] = 8'b1010100;
DRAM[12008] = 8'b1010011;
DRAM[12009] = 8'b1010100;
DRAM[12010] = 8'b1010100;
DRAM[12011] = 8'b1010101;
DRAM[12012] = 8'b1010101;
DRAM[12013] = 8'b1010100;
DRAM[12014] = 8'b1010100;
DRAM[12015] = 8'b1010011;
DRAM[12016] = 8'b1010010;
DRAM[12017] = 8'b1010010;
DRAM[12018] = 8'b1010010;
DRAM[12019] = 8'b1010001;
DRAM[12020] = 8'b1010001;
DRAM[12021] = 8'b1010000;
DRAM[12022] = 8'b1010000;
DRAM[12023] = 8'b1010000;
DRAM[12024] = 8'b1001111;
DRAM[12025] = 8'b1001111;
DRAM[12026] = 8'b1001111;
DRAM[12027] = 8'b1001111;
DRAM[12028] = 8'b1001111;
DRAM[12029] = 8'b1001111;
DRAM[12030] = 8'b1001111;
DRAM[12031] = 8'b1001111;
DRAM[12032] = 8'b1100010;
DRAM[12033] = 8'b1100010;
DRAM[12034] = 8'b1100011;
DRAM[12035] = 8'b1100100;
DRAM[12036] = 8'b1100100;
DRAM[12037] = 8'b1100101;
DRAM[12038] = 8'b1100110;
DRAM[12039] = 8'b1100110;
DRAM[12040] = 8'b1100110;
DRAM[12041] = 8'b1100110;
DRAM[12042] = 8'b1100111;
DRAM[12043] = 8'b1101000;
DRAM[12044] = 8'b1101000;
DRAM[12045] = 8'b1101001;
DRAM[12046] = 8'b1101010;
DRAM[12047] = 8'b1101010;
DRAM[12048] = 8'b1101010;
DRAM[12049] = 8'b1101010;
DRAM[12050] = 8'b1101011;
DRAM[12051] = 8'b1101100;
DRAM[12052] = 8'b1101100;
DRAM[12053] = 8'b1101101;
DRAM[12054] = 8'b1101110;
DRAM[12055] = 8'b1101110;
DRAM[12056] = 8'b1101111;
DRAM[12057] = 8'b1101110;
DRAM[12058] = 8'b1101101;
DRAM[12059] = 8'b1101101;
DRAM[12060] = 8'b1101110;
DRAM[12061] = 8'b1110000;
DRAM[12062] = 8'b1110001;
DRAM[12063] = 8'b1110011;
DRAM[12064] = 8'b1110011;
DRAM[12065] = 8'b1110011;
DRAM[12066] = 8'b1110011;
DRAM[12067] = 8'b1110100;
DRAM[12068] = 8'b1110100;
DRAM[12069] = 8'b1110101;
DRAM[12070] = 8'b1110101;
DRAM[12071] = 8'b1110101;
DRAM[12072] = 8'b1110100;
DRAM[12073] = 8'b1110100;
DRAM[12074] = 8'b1110101;
DRAM[12075] = 8'b1110110;
DRAM[12076] = 8'b1110110;
DRAM[12077] = 8'b1110111;
DRAM[12078] = 8'b1111000;
DRAM[12079] = 8'b1111000;
DRAM[12080] = 8'b1111001;
DRAM[12081] = 8'b1111001;
DRAM[12082] = 8'b1111000;
DRAM[12083] = 8'b1111010;
DRAM[12084] = 8'b1111100;
DRAM[12085] = 8'b1111100;
DRAM[12086] = 8'b1111011;
DRAM[12087] = 8'b1111001;
DRAM[12088] = 8'b1111100;
DRAM[12089] = 8'b1111011;
DRAM[12090] = 8'b1111001;
DRAM[12091] = 8'b1111000;
DRAM[12092] = 8'b1111000;
DRAM[12093] = 8'b1111010;
DRAM[12094] = 8'b1111100;
DRAM[12095] = 8'b1111110;
DRAM[12096] = 8'b10100001;
DRAM[12097] = 8'b10111100;
DRAM[12098] = 8'b11010011;
DRAM[12099] = 8'b11011001;
DRAM[12100] = 8'b11011100;
DRAM[12101] = 8'b11101000;
DRAM[12102] = 8'b11110011;
DRAM[12103] = 8'b11110111;
DRAM[12104] = 8'b11111111;
DRAM[12105] = 8'b11111010;
DRAM[12106] = 8'b11110101;
DRAM[12107] = 8'b11111110;
DRAM[12108] = 8'b11111111;
DRAM[12109] = 8'b11111000;
DRAM[12110] = 8'b11110010;
DRAM[12111] = 8'b11111111;
DRAM[12112] = 8'b11111000;
DRAM[12113] = 8'b11111111;
DRAM[12114] = 8'b11111111;
DRAM[12115] = 8'b11111111;
DRAM[12116] = 8'b11111101;
DRAM[12117] = 8'b11111101;
DRAM[12118] = 8'b11111101;
DRAM[12119] = 8'b11111011;
DRAM[12120] = 8'b11111111;
DRAM[12121] = 8'b11111111;
DRAM[12122] = 8'b11111111;
DRAM[12123] = 8'b11111111;
DRAM[12124] = 8'b11111111;
DRAM[12125] = 8'b11111111;
DRAM[12126] = 8'b11111110;
DRAM[12127] = 8'b11111101;
DRAM[12128] = 8'b11111111;
DRAM[12129] = 8'b11111111;
DRAM[12130] = 8'b11111111;
DRAM[12131] = 8'b11111111;
DRAM[12132] = 8'b11111111;
DRAM[12133] = 8'b11111111;
DRAM[12134] = 8'b11111111;
DRAM[12135] = 8'b11111111;
DRAM[12136] = 8'b11111110;
DRAM[12137] = 8'b11111110;
DRAM[12138] = 8'b11111110;
DRAM[12139] = 8'b11111110;
DRAM[12140] = 8'b11111110;
DRAM[12141] = 8'b11111110;
DRAM[12142] = 8'b11111110;
DRAM[12143] = 8'b11111110;
DRAM[12144] = 8'b11111110;
DRAM[12145] = 8'b11111110;
DRAM[12146] = 8'b11111110;
DRAM[12147] = 8'b11111110;
DRAM[12148] = 8'b11111110;
DRAM[12149] = 8'b11111110;
DRAM[12150] = 8'b11111110;
DRAM[12151] = 8'b11111110;
DRAM[12152] = 8'b11111110;
DRAM[12153] = 8'b11111110;
DRAM[12154] = 8'b11111110;
DRAM[12155] = 8'b11111111;
DRAM[12156] = 8'b11111111;
DRAM[12157] = 8'b11111111;
DRAM[12158] = 8'b11111111;
DRAM[12159] = 8'b11111111;
DRAM[12160] = 8'b11111111;
DRAM[12161] = 8'b11111111;
DRAM[12162] = 8'b11111111;
DRAM[12163] = 8'b11111111;
DRAM[12164] = 8'b11111111;
DRAM[12165] = 8'b11111111;
DRAM[12166] = 8'b11111111;
DRAM[12167] = 8'b11111111;
DRAM[12168] = 8'b11111111;
DRAM[12169] = 8'b11111111;
DRAM[12170] = 8'b11111111;
DRAM[12171] = 8'b11111111;
DRAM[12172] = 8'b11111111;
DRAM[12173] = 8'b11111111;
DRAM[12174] = 8'b11111111;
DRAM[12175] = 8'b11111111;
DRAM[12176] = 8'b11111111;
DRAM[12177] = 8'b11111111;
DRAM[12178] = 8'b11111111;
DRAM[12179] = 8'b11111110;
DRAM[12180] = 8'b11111110;
DRAM[12181] = 8'b11111101;
DRAM[12182] = 8'b11111101;
DRAM[12183] = 8'b11111101;
DRAM[12184] = 8'b11111110;
DRAM[12185] = 8'b11111110;
DRAM[12186] = 8'b11111110;
DRAM[12187] = 8'b11111111;
DRAM[12188] = 8'b11111111;
DRAM[12189] = 8'b11111111;
DRAM[12190] = 8'b11111111;
DRAM[12191] = 8'b11111111;
DRAM[12192] = 8'b11111110;
DRAM[12193] = 8'b11111110;
DRAM[12194] = 8'b11111110;
DRAM[12195] = 8'b11111110;
DRAM[12196] = 8'b11111110;
DRAM[12197] = 8'b11111110;
DRAM[12198] = 8'b11111110;
DRAM[12199] = 8'b11111110;
DRAM[12200] = 8'b11111101;
DRAM[12201] = 8'b11111101;
DRAM[12202] = 8'b11111101;
DRAM[12203] = 8'b11111110;
DRAM[12204] = 8'b11111110;
DRAM[12205] = 8'b11111111;
DRAM[12206] = 8'b11111111;
DRAM[12207] = 8'b11111111;
DRAM[12208] = 8'b11111111;
DRAM[12209] = 8'b11111111;
DRAM[12210] = 8'b11111111;
DRAM[12211] = 8'b11111111;
DRAM[12212] = 8'b11111111;
DRAM[12213] = 8'b11111111;
DRAM[12214] = 8'b11111111;
DRAM[12215] = 8'b11111111;
DRAM[12216] = 8'b11111111;
DRAM[12217] = 8'b11111111;
DRAM[12218] = 8'b11111110;
DRAM[12219] = 8'b11111111;
DRAM[12220] = 8'b11111111;
DRAM[12221] = 8'b11111100;
DRAM[12222] = 8'b11111011;
DRAM[12223] = 8'b11111100;
DRAM[12224] = 8'b11110011;
DRAM[12225] = 8'b11111111;
DRAM[12226] = 8'b11111111;
DRAM[12227] = 8'b11110110;
DRAM[12228] = 8'b11111000;
DRAM[12229] = 8'b11111011;
DRAM[12230] = 8'b11111110;
DRAM[12231] = 8'b11111111;
DRAM[12232] = 8'b11111011;
DRAM[12233] = 8'b11111011;
DRAM[12234] = 8'b11111100;
DRAM[12235] = 8'b11111001;
DRAM[12236] = 8'b11101011;
DRAM[12237] = 8'b11001100;
DRAM[12238] = 8'b10100100;
DRAM[12239] = 8'b10000111;
DRAM[12240] = 8'b1101101;
DRAM[12241] = 8'b1100110;
DRAM[12242] = 8'b1011111;
DRAM[12243] = 8'b1011101;
DRAM[12244] = 8'b1011111;
DRAM[12245] = 8'b1100010;
DRAM[12246] = 8'b1100001;
DRAM[12247] = 8'b1011111;
DRAM[12248] = 8'b1011100;
DRAM[12249] = 8'b1011100;
DRAM[12250] = 8'b1011011;
DRAM[12251] = 8'b1011010;
DRAM[12252] = 8'b1011010;
DRAM[12253] = 8'b1011001;
DRAM[12254] = 8'b1011000;
DRAM[12255] = 8'b1011000;
DRAM[12256] = 8'b1010110;
DRAM[12257] = 8'b1010110;
DRAM[12258] = 8'b1010110;
DRAM[12259] = 8'b1010101;
DRAM[12260] = 8'b1010101;
DRAM[12261] = 8'b1010100;
DRAM[12262] = 8'b1010100;
DRAM[12263] = 8'b1010100;
DRAM[12264] = 8'b1010011;
DRAM[12265] = 8'b1010100;
DRAM[12266] = 8'b1010100;
DRAM[12267] = 8'b1010101;
DRAM[12268] = 8'b1010101;
DRAM[12269] = 8'b1010100;
DRAM[12270] = 8'b1010100;
DRAM[12271] = 8'b1010011;
DRAM[12272] = 8'b1010010;
DRAM[12273] = 8'b1010010;
DRAM[12274] = 8'b1010010;
DRAM[12275] = 8'b1010001;
DRAM[12276] = 8'b1010001;
DRAM[12277] = 8'b1010000;
DRAM[12278] = 8'b1010000;
DRAM[12279] = 8'b1010000;
DRAM[12280] = 8'b1010000;
DRAM[12281] = 8'b1010000;
DRAM[12282] = 8'b1010000;
DRAM[12283] = 8'b1010000;
DRAM[12284] = 8'b1010000;
DRAM[12285] = 8'b1010000;
DRAM[12286] = 8'b1010000;
DRAM[12287] = 8'b1010000;
DRAM[12288] = 8'b1100011;
DRAM[12289] = 8'b1100011;
DRAM[12290] = 8'b1100100;
DRAM[12291] = 8'b1100101;
DRAM[12292] = 8'b1100101;
DRAM[12293] = 8'b1100110;
DRAM[12294] = 8'b1100111;
DRAM[12295] = 8'b1100111;
DRAM[12296] = 8'b1100101;
DRAM[12297] = 8'b1100110;
DRAM[12298] = 8'b1101000;
DRAM[12299] = 8'b1101010;
DRAM[12300] = 8'b1101010;
DRAM[12301] = 8'b1101001;
DRAM[12302] = 8'b1101000;
DRAM[12303] = 8'b1100111;
DRAM[12304] = 8'b1101000;
DRAM[12305] = 8'b1101001;
DRAM[12306] = 8'b1101010;
DRAM[12307] = 8'b1101011;
DRAM[12308] = 8'b1101101;
DRAM[12309] = 8'b1101110;
DRAM[12310] = 8'b1101111;
DRAM[12311] = 8'b1110000;
DRAM[12312] = 8'b1101101;
DRAM[12313] = 8'b1101110;
DRAM[12314] = 8'b1101111;
DRAM[12315] = 8'b1110000;
DRAM[12316] = 8'b1110000;
DRAM[12317] = 8'b1110000;
DRAM[12318] = 8'b1110000;
DRAM[12319] = 8'b1101111;
DRAM[12320] = 8'b1110010;
DRAM[12321] = 8'b1110010;
DRAM[12322] = 8'b1110011;
DRAM[12323] = 8'b1110100;
DRAM[12324] = 8'b1110100;
DRAM[12325] = 8'b1110101;
DRAM[12326] = 8'b1110110;
DRAM[12327] = 8'b1110110;
DRAM[12328] = 8'b1110101;
DRAM[12329] = 8'b1110101;
DRAM[12330] = 8'b1110110;
DRAM[12331] = 8'b1110111;
DRAM[12332] = 8'b1110111;
DRAM[12333] = 8'b1111000;
DRAM[12334] = 8'b1111001;
DRAM[12335] = 8'b1111001;
DRAM[12336] = 8'b1111110;
DRAM[12337] = 8'b1110111;
DRAM[12338] = 8'b1110100;
DRAM[12339] = 8'b1111001;
DRAM[12340] = 8'b1111010;
DRAM[12341] = 8'b1111000;
DRAM[12342] = 8'b1111010;
DRAM[12343] = 8'b10000001;
DRAM[12344] = 8'b1111110;
DRAM[12345] = 8'b1111110;
DRAM[12346] = 8'b1111111;
DRAM[12347] = 8'b10000001;
DRAM[12348] = 8'b10000010;
DRAM[12349] = 8'b10000011;
DRAM[12350] = 8'b10001000;
DRAM[12351] = 8'b10001101;
DRAM[12352] = 8'b10101101;
DRAM[12353] = 8'b11001110;
DRAM[12354] = 8'b11101101;
DRAM[12355] = 8'b11110110;
DRAM[12356] = 8'b11110111;
DRAM[12357] = 8'b11111100;
DRAM[12358] = 8'b11111111;
DRAM[12359] = 8'b11111111;
DRAM[12360] = 8'b11111101;
DRAM[12361] = 8'b11111101;
DRAM[12362] = 8'b11111101;
DRAM[12363] = 8'b11111110;
DRAM[12364] = 8'b11111110;
DRAM[12365] = 8'b11111111;
DRAM[12366] = 8'b11111111;
DRAM[12367] = 8'b11111111;
DRAM[12368] = 8'b11111111;
DRAM[12369] = 8'b11111111;
DRAM[12370] = 8'b11111111;
DRAM[12371] = 8'b11111111;
DRAM[12372] = 8'b11111111;
DRAM[12373] = 8'b11111111;
DRAM[12374] = 8'b11111111;
DRAM[12375] = 8'b11111111;
DRAM[12376] = 8'b11111111;
DRAM[12377] = 8'b11111111;
DRAM[12378] = 8'b11111111;
DRAM[12379] = 8'b11111111;
DRAM[12380] = 8'b11111111;
DRAM[12381] = 8'b11111111;
DRAM[12382] = 8'b11111111;
DRAM[12383] = 8'b11111111;
DRAM[12384] = 8'b11111101;
DRAM[12385] = 8'b11111110;
DRAM[12386] = 8'b11111110;
DRAM[12387] = 8'b11111110;
DRAM[12388] = 8'b11111110;
DRAM[12389] = 8'b11111101;
DRAM[12390] = 8'b11111100;
DRAM[12391] = 8'b11111011;
DRAM[12392] = 8'b11111111;
DRAM[12393] = 8'b11111111;
DRAM[12394] = 8'b11111111;
DRAM[12395] = 8'b11111111;
DRAM[12396] = 8'b11111110;
DRAM[12397] = 8'b11111101;
DRAM[12398] = 8'b11111100;
DRAM[12399] = 8'b11111011;
DRAM[12400] = 8'b11111111;
DRAM[12401] = 8'b11111111;
DRAM[12402] = 8'b11111110;
DRAM[12403] = 8'b11111101;
DRAM[12404] = 8'b11111101;
DRAM[12405] = 8'b11111110;
DRAM[12406] = 8'b11111110;
DRAM[12407] = 8'b11111110;
DRAM[12408] = 8'b11111110;
DRAM[12409] = 8'b11111110;
DRAM[12410] = 8'b11111111;
DRAM[12411] = 8'b11111111;
DRAM[12412] = 8'b11111111;
DRAM[12413] = 8'b11111111;
DRAM[12414] = 8'b11111111;
DRAM[12415] = 8'b11111111;
DRAM[12416] = 8'b11111111;
DRAM[12417] = 8'b11111111;
DRAM[12418] = 8'b11111110;
DRAM[12419] = 8'b11111101;
DRAM[12420] = 8'b11111110;
DRAM[12421] = 8'b11111111;
DRAM[12422] = 8'b11111111;
DRAM[12423] = 8'b11111111;
DRAM[12424] = 8'b11111100;
DRAM[12425] = 8'b11111100;
DRAM[12426] = 8'b11111101;
DRAM[12427] = 8'b11111110;
DRAM[12428] = 8'b11111110;
DRAM[12429] = 8'b11111101;
DRAM[12430] = 8'b11111101;
DRAM[12431] = 8'b11111100;
DRAM[12432] = 8'b11111100;
DRAM[12433] = 8'b11111101;
DRAM[12434] = 8'b11111101;
DRAM[12435] = 8'b11111101;
DRAM[12436] = 8'b11111101;
DRAM[12437] = 8'b11111100;
DRAM[12438] = 8'b11111011;
DRAM[12439] = 8'b11111010;
DRAM[12440] = 8'b11111011;
DRAM[12441] = 8'b11111011;
DRAM[12442] = 8'b11111100;
DRAM[12443] = 8'b11111100;
DRAM[12444] = 8'b11111100;
DRAM[12445] = 8'b11111100;
DRAM[12446] = 8'b11111101;
DRAM[12447] = 8'b11111101;
DRAM[12448] = 8'b11111111;
DRAM[12449] = 8'b11111111;
DRAM[12450] = 8'b11111111;
DRAM[12451] = 8'b11111111;
DRAM[12452] = 8'b11111111;
DRAM[12453] = 8'b11111111;
DRAM[12454] = 8'b11111111;
DRAM[12455] = 8'b11111111;
DRAM[12456] = 8'b11111100;
DRAM[12457] = 8'b11111100;
DRAM[12458] = 8'b11111100;
DRAM[12459] = 8'b11111101;
DRAM[12460] = 8'b11111101;
DRAM[12461] = 8'b11111110;
DRAM[12462] = 8'b11111110;
DRAM[12463] = 8'b11111110;
DRAM[12464] = 8'b11111111;
DRAM[12465] = 8'b11111111;
DRAM[12466] = 8'b11111111;
DRAM[12467] = 8'b11111101;
DRAM[12468] = 8'b11111100;
DRAM[12469] = 8'b11111011;
DRAM[12470] = 8'b11111011;
DRAM[12471] = 8'b11111011;
DRAM[12472] = 8'b11111100;
DRAM[12473] = 8'b11111101;
DRAM[12474] = 8'b11111111;
DRAM[12475] = 8'b11111110;
DRAM[12476] = 8'b11111101;
DRAM[12477] = 8'b11111011;
DRAM[12478] = 8'b11111010;
DRAM[12479] = 8'b11111010;
DRAM[12480] = 8'b11111110;
DRAM[12481] = 8'b11111110;
DRAM[12482] = 8'b11111110;
DRAM[12483] = 8'b11111110;
DRAM[12484] = 8'b11111110;
DRAM[12485] = 8'b11111110;
DRAM[12486] = 8'b11111110;
DRAM[12487] = 8'b11111110;
DRAM[12488] = 8'b11111100;
DRAM[12489] = 8'b11111100;
DRAM[12490] = 8'b11111011;
DRAM[12491] = 8'b11111100;
DRAM[12492] = 8'b11111101;
DRAM[12493] = 8'b11101011;
DRAM[12494] = 8'b10111011;
DRAM[12495] = 8'b10001011;
DRAM[12496] = 8'b10001110;
DRAM[12497] = 8'b10010100;
DRAM[12498] = 8'b10100001;
DRAM[12499] = 8'b10011101;
DRAM[12500] = 8'b10001000;
DRAM[12501] = 8'b1111100;
DRAM[12502] = 8'b1110110;
DRAM[12503] = 8'b1101011;
DRAM[12504] = 8'b1101001;
DRAM[12505] = 8'b1100010;
DRAM[12506] = 8'b1011110;
DRAM[12507] = 8'b1011101;
DRAM[12508] = 8'b1011011;
DRAM[12509] = 8'b1011001;
DRAM[12510] = 8'b1011010;
DRAM[12511] = 8'b1011110;
DRAM[12512] = 8'b1010111;
DRAM[12513] = 8'b1010111;
DRAM[12514] = 8'b1010111;
DRAM[12515] = 8'b1010110;
DRAM[12516] = 8'b1010110;
DRAM[12517] = 8'b1010101;
DRAM[12518] = 8'b1010101;
DRAM[12519] = 8'b1010101;
DRAM[12520] = 8'b1010100;
DRAM[12521] = 8'b1010100;
DRAM[12522] = 8'b1010011;
DRAM[12523] = 8'b1010011;
DRAM[12524] = 8'b1010011;
DRAM[12525] = 8'b1010010;
DRAM[12526] = 8'b1010010;
DRAM[12527] = 8'b1010010;
DRAM[12528] = 8'b1010010;
DRAM[12529] = 8'b1010010;
DRAM[12530] = 8'b1010010;
DRAM[12531] = 8'b1010001;
DRAM[12532] = 8'b1010001;
DRAM[12533] = 8'b1010000;
DRAM[12534] = 8'b1010000;
DRAM[12535] = 8'b1010000;
DRAM[12536] = 8'b1010000;
DRAM[12537] = 8'b1010000;
DRAM[12538] = 8'b1010000;
DRAM[12539] = 8'b1010000;
DRAM[12540] = 8'b1010000;
DRAM[12541] = 8'b1010000;
DRAM[12542] = 8'b1010000;
DRAM[12543] = 8'b1010000;
DRAM[12544] = 8'b1100011;
DRAM[12545] = 8'b1100011;
DRAM[12546] = 8'b1100100;
DRAM[12547] = 8'b1100101;
DRAM[12548] = 8'b1100101;
DRAM[12549] = 8'b1100110;
DRAM[12550] = 8'b1100111;
DRAM[12551] = 8'b1100111;
DRAM[12552] = 8'b1100110;
DRAM[12553] = 8'b1100111;
DRAM[12554] = 8'b1101000;
DRAM[12555] = 8'b1101000;
DRAM[12556] = 8'b1101001;
DRAM[12557] = 8'b1101001;
DRAM[12558] = 8'b1101001;
DRAM[12559] = 8'b1101000;
DRAM[12560] = 8'b1101001;
DRAM[12561] = 8'b1101010;
DRAM[12562] = 8'b1101010;
DRAM[12563] = 8'b1101011;
DRAM[12564] = 8'b1101101;
DRAM[12565] = 8'b1101110;
DRAM[12566] = 8'b1101110;
DRAM[12567] = 8'b1101111;
DRAM[12568] = 8'b1101101;
DRAM[12569] = 8'b1101110;
DRAM[12570] = 8'b1101111;
DRAM[12571] = 8'b1110000;
DRAM[12572] = 8'b1110000;
DRAM[12573] = 8'b1110000;
DRAM[12574] = 8'b1110000;
DRAM[12575] = 8'b1101111;
DRAM[12576] = 8'b1110010;
DRAM[12577] = 8'b1110010;
DRAM[12578] = 8'b1110011;
DRAM[12579] = 8'b1110100;
DRAM[12580] = 8'b1110100;
DRAM[12581] = 8'b1110101;
DRAM[12582] = 8'b1110110;
DRAM[12583] = 8'b1110110;
DRAM[12584] = 8'b1110101;
DRAM[12585] = 8'b1110101;
DRAM[12586] = 8'b1110110;
DRAM[12587] = 8'b1110111;
DRAM[12588] = 8'b1111000;
DRAM[12589] = 8'b1111000;
DRAM[12590] = 8'b1111001;
DRAM[12591] = 8'b1111001;
DRAM[12592] = 8'b1110111;
DRAM[12593] = 8'b1111000;
DRAM[12594] = 8'b1111100;
DRAM[12595] = 8'b10000000;
DRAM[12596] = 8'b10000001;
DRAM[12597] = 8'b1111111;
DRAM[12598] = 8'b1111111;
DRAM[12599] = 8'b10000001;
DRAM[12600] = 8'b10000100;
DRAM[12601] = 8'b10000001;
DRAM[12602] = 8'b1111110;
DRAM[12603] = 8'b1111101;
DRAM[12604] = 8'b10000001;
DRAM[12605] = 8'b10001101;
DRAM[12606] = 8'b10011110;
DRAM[12607] = 8'b10101011;
DRAM[12608] = 8'b11000001;
DRAM[12609] = 8'b11011011;
DRAM[12610] = 8'b11110011;
DRAM[12611] = 8'b11111001;
DRAM[12612] = 8'b11111010;
DRAM[12613] = 8'b11111110;
DRAM[12614] = 8'b11111111;
DRAM[12615] = 8'b11111110;
DRAM[12616] = 8'b11111101;
DRAM[12617] = 8'b11111101;
DRAM[12618] = 8'b11111101;
DRAM[12619] = 8'b11111110;
DRAM[12620] = 8'b11111110;
DRAM[12621] = 8'b11111111;
DRAM[12622] = 8'b11111111;
DRAM[12623] = 8'b11111111;
DRAM[12624] = 8'b11111111;
DRAM[12625] = 8'b11111111;
DRAM[12626] = 8'b11111111;
DRAM[12627] = 8'b11111111;
DRAM[12628] = 8'b11111111;
DRAM[12629] = 8'b11111111;
DRAM[12630] = 8'b11111111;
DRAM[12631] = 8'b11111111;
DRAM[12632] = 8'b11111111;
DRAM[12633] = 8'b11111111;
DRAM[12634] = 8'b11111111;
DRAM[12635] = 8'b11111111;
DRAM[12636] = 8'b11111111;
DRAM[12637] = 8'b11111111;
DRAM[12638] = 8'b11111111;
DRAM[12639] = 8'b11111111;
DRAM[12640] = 8'b11111101;
DRAM[12641] = 8'b11111110;
DRAM[12642] = 8'b11111110;
DRAM[12643] = 8'b11111110;
DRAM[12644] = 8'b11111110;
DRAM[12645] = 8'b11111101;
DRAM[12646] = 8'b11111100;
DRAM[12647] = 8'b11111011;
DRAM[12648] = 8'b11111111;
DRAM[12649] = 8'b11111111;
DRAM[12650] = 8'b11111111;
DRAM[12651] = 8'b11111111;
DRAM[12652] = 8'b11111110;
DRAM[12653] = 8'b11111101;
DRAM[12654] = 8'b11111100;
DRAM[12655] = 8'b11111011;
DRAM[12656] = 8'b11111110;
DRAM[12657] = 8'b11111110;
DRAM[12658] = 8'b11111110;
DRAM[12659] = 8'b11111101;
DRAM[12660] = 8'b11111101;
DRAM[12661] = 8'b11111101;
DRAM[12662] = 8'b11111110;
DRAM[12663] = 8'b11111110;
DRAM[12664] = 8'b11111100;
DRAM[12665] = 8'b11111101;
DRAM[12666] = 8'b11111101;
DRAM[12667] = 8'b11111101;
DRAM[12668] = 8'b11111110;
DRAM[12669] = 8'b11111110;
DRAM[12670] = 8'b11111110;
DRAM[12671] = 8'b11111111;
DRAM[12672] = 8'b11111110;
DRAM[12673] = 8'b11111110;
DRAM[12674] = 8'b11111101;
DRAM[12675] = 8'b11111101;
DRAM[12676] = 8'b11111101;
DRAM[12677] = 8'b11111110;
DRAM[12678] = 8'b11111111;
DRAM[12679] = 8'b11111111;
DRAM[12680] = 8'b11111100;
DRAM[12681] = 8'b11111101;
DRAM[12682] = 8'b11111110;
DRAM[12683] = 8'b11111110;
DRAM[12684] = 8'b11111110;
DRAM[12685] = 8'b11111110;
DRAM[12686] = 8'b11111101;
DRAM[12687] = 8'b11111101;
DRAM[12688] = 8'b11111101;
DRAM[12689] = 8'b11111101;
DRAM[12690] = 8'b11111101;
DRAM[12691] = 8'b11111101;
DRAM[12692] = 8'b11111100;
DRAM[12693] = 8'b11111100;
DRAM[12694] = 8'b11111011;
DRAM[12695] = 8'b11111010;
DRAM[12696] = 8'b11111011;
DRAM[12697] = 8'b11111011;
DRAM[12698] = 8'b11111100;
DRAM[12699] = 8'b11111100;
DRAM[12700] = 8'b11111100;
DRAM[12701] = 8'b11111101;
DRAM[12702] = 8'b11111101;
DRAM[12703] = 8'b11111101;
DRAM[12704] = 8'b11111111;
DRAM[12705] = 8'b11111111;
DRAM[12706] = 8'b11111111;
DRAM[12707] = 8'b11111111;
DRAM[12708] = 8'b11111111;
DRAM[12709] = 8'b11111111;
DRAM[12710] = 8'b11111111;
DRAM[12711] = 8'b11111111;
DRAM[12712] = 8'b11111101;
DRAM[12713] = 8'b11111101;
DRAM[12714] = 8'b11111101;
DRAM[12715] = 8'b11111110;
DRAM[12716] = 8'b11111110;
DRAM[12717] = 8'b11111111;
DRAM[12718] = 8'b11111111;
DRAM[12719] = 8'b11111111;
DRAM[12720] = 8'b11111111;
DRAM[12721] = 8'b11111110;
DRAM[12722] = 8'b11111011;
DRAM[12723] = 8'b11111011;
DRAM[12724] = 8'b11111101;
DRAM[12725] = 8'b11111110;
DRAM[12726] = 8'b11111110;
DRAM[12727] = 8'b11111100;
DRAM[12728] = 8'b11111011;
DRAM[12729] = 8'b11111101;
DRAM[12730] = 8'b11111110;
DRAM[12731] = 8'b11111110;
DRAM[12732] = 8'b11111100;
DRAM[12733] = 8'b11111100;
DRAM[12734] = 8'b11111110;
DRAM[12735] = 8'b11111111;
DRAM[12736] = 8'b11111110;
DRAM[12737] = 8'b11111110;
DRAM[12738] = 8'b11111110;
DRAM[12739] = 8'b11111110;
DRAM[12740] = 8'b11111110;
DRAM[12741] = 8'b11111110;
DRAM[12742] = 8'b11111110;
DRAM[12743] = 8'b11111110;
DRAM[12744] = 8'b11111110;
DRAM[12745] = 8'b11111111;
DRAM[12746] = 8'b11111100;
DRAM[12747] = 8'b11111000;
DRAM[12748] = 8'b11111000;
DRAM[12749] = 8'b11110100;
DRAM[12750] = 8'b11011101;
DRAM[12751] = 8'b11000100;
DRAM[12752] = 8'b11010011;
DRAM[12753] = 8'b10111100;
DRAM[12754] = 8'b10101001;
DRAM[12755] = 8'b10011010;
DRAM[12756] = 8'b10001010;
DRAM[12757] = 8'b10000010;
DRAM[12758] = 8'b1111011;
DRAM[12759] = 8'b1101110;
DRAM[12760] = 8'b1101000;
DRAM[12761] = 8'b1100010;
DRAM[12762] = 8'b1011110;
DRAM[12763] = 8'b1011110;
DRAM[12764] = 8'b1011100;
DRAM[12765] = 8'b1011001;
DRAM[12766] = 8'b1011001;
DRAM[12767] = 8'b1011011;
DRAM[12768] = 8'b1010111;
DRAM[12769] = 8'b1010111;
DRAM[12770] = 8'b1010111;
DRAM[12771] = 8'b1010110;
DRAM[12772] = 8'b1010110;
DRAM[12773] = 8'b1010110;
DRAM[12774] = 8'b1010101;
DRAM[12775] = 8'b1010101;
DRAM[12776] = 8'b1010110;
DRAM[12777] = 8'b1010110;
DRAM[12778] = 8'b1010110;
DRAM[12779] = 8'b1010101;
DRAM[12780] = 8'b1010101;
DRAM[12781] = 8'b1010101;
DRAM[12782] = 8'b1010100;
DRAM[12783] = 8'b1010100;
DRAM[12784] = 8'b1010010;
DRAM[12785] = 8'b1010010;
DRAM[12786] = 8'b1010010;
DRAM[12787] = 8'b1010001;
DRAM[12788] = 8'b1010001;
DRAM[12789] = 8'b1010001;
DRAM[12790] = 8'b1010000;
DRAM[12791] = 8'b1010000;
DRAM[12792] = 8'b1010000;
DRAM[12793] = 8'b1010000;
DRAM[12794] = 8'b1010000;
DRAM[12795] = 8'b1010000;
DRAM[12796] = 8'b1010000;
DRAM[12797] = 8'b1010000;
DRAM[12798] = 8'b1010000;
DRAM[12799] = 8'b1010000;
DRAM[12800] = 8'b1100011;
DRAM[12801] = 8'b1100011;
DRAM[12802] = 8'b1100100;
DRAM[12803] = 8'b1100101;
DRAM[12804] = 8'b1100101;
DRAM[12805] = 8'b1100110;
DRAM[12806] = 8'b1100111;
DRAM[12807] = 8'b1100111;
DRAM[12808] = 8'b1101000;
DRAM[12809] = 8'b1100111;
DRAM[12810] = 8'b1100111;
DRAM[12811] = 8'b1100111;
DRAM[12812] = 8'b1101000;
DRAM[12813] = 8'b1101000;
DRAM[12814] = 8'b1101001;
DRAM[12815] = 8'b1101010;
DRAM[12816] = 8'b1101011;
DRAM[12817] = 8'b1101011;
DRAM[12818] = 8'b1101011;
DRAM[12819] = 8'b1101100;
DRAM[12820] = 8'b1101100;
DRAM[12821] = 8'b1101101;
DRAM[12822] = 8'b1101101;
DRAM[12823] = 8'b1101101;
DRAM[12824] = 8'b1101101;
DRAM[12825] = 8'b1101110;
DRAM[12826] = 8'b1101111;
DRAM[12827] = 8'b1110000;
DRAM[12828] = 8'b1110000;
DRAM[12829] = 8'b1110000;
DRAM[12830] = 8'b1110000;
DRAM[12831] = 8'b1101111;
DRAM[12832] = 8'b1110010;
DRAM[12833] = 8'b1110010;
DRAM[12834] = 8'b1110011;
DRAM[12835] = 8'b1110100;
DRAM[12836] = 8'b1110100;
DRAM[12837] = 8'b1110101;
DRAM[12838] = 8'b1110110;
DRAM[12839] = 8'b1110110;
DRAM[12840] = 8'b1110101;
DRAM[12841] = 8'b1110110;
DRAM[12842] = 8'b1110110;
DRAM[12843] = 8'b1110111;
DRAM[12844] = 8'b1111000;
DRAM[12845] = 8'b1111001;
DRAM[12846] = 8'b1111001;
DRAM[12847] = 8'b1111001;
DRAM[12848] = 8'b1110111;
DRAM[12849] = 8'b1111100;
DRAM[12850] = 8'b10000000;
DRAM[12851] = 8'b1111111;
DRAM[12852] = 8'b1111101;
DRAM[12853] = 8'b1111110;
DRAM[12854] = 8'b1111110;
DRAM[12855] = 8'b1111100;
DRAM[12856] = 8'b1111101;
DRAM[12857] = 8'b10000001;
DRAM[12858] = 8'b10000101;
DRAM[12859] = 8'b10000111;
DRAM[12860] = 8'b10001010;
DRAM[12861] = 8'b10010010;
DRAM[12862] = 8'b10011100;
DRAM[12863] = 8'b10100011;
DRAM[12864] = 8'b11011100;
DRAM[12865] = 8'b11101101;
DRAM[12866] = 8'b11111010;
DRAM[12867] = 8'b11111100;
DRAM[12868] = 8'b11111100;
DRAM[12869] = 8'b11111111;
DRAM[12870] = 8'b11111111;
DRAM[12871] = 8'b11111101;
DRAM[12872] = 8'b11111101;
DRAM[12873] = 8'b11111101;
DRAM[12874] = 8'b11111110;
DRAM[12875] = 8'b11111110;
DRAM[12876] = 8'b11111110;
DRAM[12877] = 8'b11111110;
DRAM[12878] = 8'b11111111;
DRAM[12879] = 8'b11111111;
DRAM[12880] = 8'b11111111;
DRAM[12881] = 8'b11111111;
DRAM[12882] = 8'b11111111;
DRAM[12883] = 8'b11111111;
DRAM[12884] = 8'b11111111;
DRAM[12885] = 8'b11111111;
DRAM[12886] = 8'b11111111;
DRAM[12887] = 8'b11111111;
DRAM[12888] = 8'b11111111;
DRAM[12889] = 8'b11111111;
DRAM[12890] = 8'b11111111;
DRAM[12891] = 8'b11111111;
DRAM[12892] = 8'b11111111;
DRAM[12893] = 8'b11111111;
DRAM[12894] = 8'b11111111;
DRAM[12895] = 8'b11111111;
DRAM[12896] = 8'b11111101;
DRAM[12897] = 8'b11111110;
DRAM[12898] = 8'b11111110;
DRAM[12899] = 8'b11111110;
DRAM[12900] = 8'b11111110;
DRAM[12901] = 8'b11111101;
DRAM[12902] = 8'b11111100;
DRAM[12903] = 8'b11111011;
DRAM[12904] = 8'b11111101;
DRAM[12905] = 8'b11111101;
DRAM[12906] = 8'b11111110;
DRAM[12907] = 8'b11111110;
DRAM[12908] = 8'b11111110;
DRAM[12909] = 8'b11111101;
DRAM[12910] = 8'b11111101;
DRAM[12911] = 8'b11111100;
DRAM[12912] = 8'b11111101;
DRAM[12913] = 8'b11111101;
DRAM[12914] = 8'b11111101;
DRAM[12915] = 8'b11111101;
DRAM[12916] = 8'b11111101;
DRAM[12917] = 8'b11111101;
DRAM[12918] = 8'b11111101;
DRAM[12919] = 8'b11111101;
DRAM[12920] = 8'b11111011;
DRAM[12921] = 8'b11111011;
DRAM[12922] = 8'b11111011;
DRAM[12923] = 8'b11111100;
DRAM[12924] = 8'b11111100;
DRAM[12925] = 8'b11111101;
DRAM[12926] = 8'b11111101;
DRAM[12927] = 8'b11111101;
DRAM[12928] = 8'b11111110;
DRAM[12929] = 8'b11111101;
DRAM[12930] = 8'b11111101;
DRAM[12931] = 8'b11111101;
DRAM[12932] = 8'b11111101;
DRAM[12933] = 8'b11111110;
DRAM[12934] = 8'b11111111;
DRAM[12935] = 8'b11111111;
DRAM[12936] = 8'b11111101;
DRAM[12937] = 8'b11111110;
DRAM[12938] = 8'b11111111;
DRAM[12939] = 8'b11111111;
DRAM[12940] = 8'b11111111;
DRAM[12941] = 8'b11111110;
DRAM[12942] = 8'b11111110;
DRAM[12943] = 8'b11111101;
DRAM[12944] = 8'b11111101;
DRAM[12945] = 8'b11111101;
DRAM[12946] = 8'b11111100;
DRAM[12947] = 8'b11111100;
DRAM[12948] = 8'b11111100;
DRAM[12949] = 8'b11111011;
DRAM[12950] = 8'b11111011;
DRAM[12951] = 8'b11111011;
DRAM[12952] = 8'b11111011;
DRAM[12953] = 8'b11111011;
DRAM[12954] = 8'b11111100;
DRAM[12955] = 8'b11111100;
DRAM[12956] = 8'b11111101;
DRAM[12957] = 8'b11111101;
DRAM[12958] = 8'b11111101;
DRAM[12959] = 8'b11111110;
DRAM[12960] = 8'b11111111;
DRAM[12961] = 8'b11111111;
DRAM[12962] = 8'b11111111;
DRAM[12963] = 8'b11111111;
DRAM[12964] = 8'b11111111;
DRAM[12965] = 8'b11111111;
DRAM[12966] = 8'b11111111;
DRAM[12967] = 8'b11111111;
DRAM[12968] = 8'b11111110;
DRAM[12969] = 8'b11111110;
DRAM[12970] = 8'b11111110;
DRAM[12971] = 8'b11111111;
DRAM[12972] = 8'b11111111;
DRAM[12973] = 8'b11111111;
DRAM[12974] = 8'b11111111;
DRAM[12975] = 8'b11111111;
DRAM[12976] = 8'b11111111;
DRAM[12977] = 8'b11111100;
DRAM[12978] = 8'b11111000;
DRAM[12979] = 8'b11111001;
DRAM[12980] = 8'b11111100;
DRAM[12981] = 8'b11111110;
DRAM[12982] = 8'b11111110;
DRAM[12983] = 8'b11111101;
DRAM[12984] = 8'b11111010;
DRAM[12985] = 8'b11111100;
DRAM[12986] = 8'b11111110;
DRAM[12987] = 8'b11111101;
DRAM[12988] = 8'b11111011;
DRAM[12989] = 8'b11111100;
DRAM[12990] = 8'b11111111;
DRAM[12991] = 8'b11111111;
DRAM[12992] = 8'b11111110;
DRAM[12993] = 8'b11111110;
DRAM[12994] = 8'b11111110;
DRAM[12995] = 8'b11111110;
DRAM[12996] = 8'b11111110;
DRAM[12997] = 8'b11111110;
DRAM[12998] = 8'b11111110;
DRAM[12999] = 8'b11111110;
DRAM[13000] = 8'b11111100;
DRAM[13001] = 8'b11111111;
DRAM[13002] = 8'b11111111;
DRAM[13003] = 8'b11111000;
DRAM[13004] = 8'b11110111;
DRAM[13005] = 8'b11111011;
DRAM[13006] = 8'b11111011;
DRAM[13007] = 8'b11110110;
DRAM[13008] = 8'b11100110;
DRAM[13009] = 8'b11000000;
DRAM[13010] = 8'b10100000;
DRAM[13011] = 8'b10001010;
DRAM[13012] = 8'b1110101;
DRAM[13013] = 8'b1101001;
DRAM[13014] = 8'b1100101;
DRAM[13015] = 8'b1011110;
DRAM[13016] = 8'b1100111;
DRAM[13017] = 8'b1100001;
DRAM[13018] = 8'b1011101;
DRAM[13019] = 8'b1011101;
DRAM[13020] = 8'b1011101;
DRAM[13021] = 8'b1011001;
DRAM[13022] = 8'b1011000;
DRAM[13023] = 8'b1011001;
DRAM[13024] = 8'b1010111;
DRAM[13025] = 8'b1010111;
DRAM[13026] = 8'b1010111;
DRAM[13027] = 8'b1010111;
DRAM[13028] = 8'b1010110;
DRAM[13029] = 8'b1010110;
DRAM[13030] = 8'b1010110;
DRAM[13031] = 8'b1010101;
DRAM[13032] = 8'b1010111;
DRAM[13033] = 8'b1010110;
DRAM[13034] = 8'b1010110;
DRAM[13035] = 8'b1010110;
DRAM[13036] = 8'b1010101;
DRAM[13037] = 8'b1010101;
DRAM[13038] = 8'b1010101;
DRAM[13039] = 8'b1010100;
DRAM[13040] = 8'b1010010;
DRAM[13041] = 8'b1010010;
DRAM[13042] = 8'b1010010;
DRAM[13043] = 8'b1010010;
DRAM[13044] = 8'b1010001;
DRAM[13045] = 8'b1010001;
DRAM[13046] = 8'b1010001;
DRAM[13047] = 8'b1010000;
DRAM[13048] = 8'b1010000;
DRAM[13049] = 8'b1010000;
DRAM[13050] = 8'b1010000;
DRAM[13051] = 8'b1010000;
DRAM[13052] = 8'b1010000;
DRAM[13053] = 8'b1010000;
DRAM[13054] = 8'b1010000;
DRAM[13055] = 8'b1010000;
DRAM[13056] = 8'b1100011;
DRAM[13057] = 8'b1100011;
DRAM[13058] = 8'b1100100;
DRAM[13059] = 8'b1100101;
DRAM[13060] = 8'b1100101;
DRAM[13061] = 8'b1100110;
DRAM[13062] = 8'b1100111;
DRAM[13063] = 8'b1100111;
DRAM[13064] = 8'b1101001;
DRAM[13065] = 8'b1101000;
DRAM[13066] = 8'b1100111;
DRAM[13067] = 8'b1100110;
DRAM[13068] = 8'b1100110;
DRAM[13069] = 8'b1101000;
DRAM[13070] = 8'b1101010;
DRAM[13071] = 8'b1101011;
DRAM[13072] = 8'b1101100;
DRAM[13073] = 8'b1101100;
DRAM[13074] = 8'b1101100;
DRAM[13075] = 8'b1101100;
DRAM[13076] = 8'b1101100;
DRAM[13077] = 8'b1101100;
DRAM[13078] = 8'b1101100;
DRAM[13079] = 8'b1101100;
DRAM[13080] = 8'b1101101;
DRAM[13081] = 8'b1101110;
DRAM[13082] = 8'b1101111;
DRAM[13083] = 8'b1110000;
DRAM[13084] = 8'b1110000;
DRAM[13085] = 8'b1110000;
DRAM[13086] = 8'b1110000;
DRAM[13087] = 8'b1101111;
DRAM[13088] = 8'b1110010;
DRAM[13089] = 8'b1110010;
DRAM[13090] = 8'b1110011;
DRAM[13091] = 8'b1110100;
DRAM[13092] = 8'b1110100;
DRAM[13093] = 8'b1110101;
DRAM[13094] = 8'b1110110;
DRAM[13095] = 8'b1110110;
DRAM[13096] = 8'b1110110;
DRAM[13097] = 8'b1110110;
DRAM[13098] = 8'b1110111;
DRAM[13099] = 8'b1110111;
DRAM[13100] = 8'b1111000;
DRAM[13101] = 8'b1111001;
DRAM[13102] = 8'b1111010;
DRAM[13103] = 8'b1111010;
DRAM[13104] = 8'b1111010;
DRAM[13105] = 8'b1111101;
DRAM[13106] = 8'b1111011;
DRAM[13107] = 8'b1111000;
DRAM[13108] = 8'b1111010;
DRAM[13109] = 8'b10000011;
DRAM[13110] = 8'b10000110;
DRAM[13111] = 8'b10000011;
DRAM[13112] = 8'b10011000;
DRAM[13113] = 8'b10010110;
DRAM[13114] = 8'b10010000;
DRAM[13115] = 8'b10001100;
DRAM[13116] = 8'b10010101;
DRAM[13117] = 8'b10101110;
DRAM[13118] = 8'b11001101;
DRAM[13119] = 8'b11100001;
DRAM[13120] = 8'b11110001;
DRAM[13121] = 8'b11111000;
DRAM[13122] = 8'b11111101;
DRAM[13123] = 8'b11111100;
DRAM[13124] = 8'b11111101;
DRAM[13125] = 8'b11111111;
DRAM[13126] = 8'b11111111;
DRAM[13127] = 8'b11111100;
DRAM[13128] = 8'b11111110;
DRAM[13129] = 8'b11111110;
DRAM[13130] = 8'b11111110;
DRAM[13131] = 8'b11111110;
DRAM[13132] = 8'b11111110;
DRAM[13133] = 8'b11111110;
DRAM[13134] = 8'b11111110;
DRAM[13135] = 8'b11111110;
DRAM[13136] = 8'b11111110;
DRAM[13137] = 8'b11111110;
DRAM[13138] = 8'b11111110;
DRAM[13139] = 8'b11111110;
DRAM[13140] = 8'b11111110;
DRAM[13141] = 8'b11111110;
DRAM[13142] = 8'b11111110;
DRAM[13143] = 8'b11111110;
DRAM[13144] = 8'b11111110;
DRAM[13145] = 8'b11111110;
DRAM[13146] = 8'b11111110;
DRAM[13147] = 8'b11111110;
DRAM[13148] = 8'b11111110;
DRAM[13149] = 8'b11111110;
DRAM[13150] = 8'b11111110;
DRAM[13151] = 8'b11111110;
DRAM[13152] = 8'b11111101;
DRAM[13153] = 8'b11111110;
DRAM[13154] = 8'b11111110;
DRAM[13155] = 8'b11111110;
DRAM[13156] = 8'b11111110;
DRAM[13157] = 8'b11111101;
DRAM[13158] = 8'b11111100;
DRAM[13159] = 8'b11111011;
DRAM[13160] = 8'b11111011;
DRAM[13161] = 8'b11111100;
DRAM[13162] = 8'b11111100;
DRAM[13163] = 8'b11111101;
DRAM[13164] = 8'b11111101;
DRAM[13165] = 8'b11111101;
DRAM[13166] = 8'b11111101;
DRAM[13167] = 8'b11111100;
DRAM[13168] = 8'b11111011;
DRAM[13169] = 8'b11111100;
DRAM[13170] = 8'b11111100;
DRAM[13171] = 8'b11111101;
DRAM[13172] = 8'b11111101;
DRAM[13173] = 8'b11111101;
DRAM[13174] = 8'b11111101;
DRAM[13175] = 8'b11111101;
DRAM[13176] = 8'b11111011;
DRAM[13177] = 8'b11111011;
DRAM[13178] = 8'b11111011;
DRAM[13179] = 8'b11111100;
DRAM[13180] = 8'b11111100;
DRAM[13181] = 8'b11111100;
DRAM[13182] = 8'b11111101;
DRAM[13183] = 8'b11111101;
DRAM[13184] = 8'b11111110;
DRAM[13185] = 8'b11111110;
DRAM[13186] = 8'b11111110;
DRAM[13187] = 8'b11111110;
DRAM[13188] = 8'b11111111;
DRAM[13189] = 8'b11111111;
DRAM[13190] = 8'b11111111;
DRAM[13191] = 8'b11111111;
DRAM[13192] = 8'b11111110;
DRAM[13193] = 8'b11111111;
DRAM[13194] = 8'b11111111;
DRAM[13195] = 8'b11111111;
DRAM[13196] = 8'b11111111;
DRAM[13197] = 8'b11111110;
DRAM[13198] = 8'b11111101;
DRAM[13199] = 8'b11111101;
DRAM[13200] = 8'b11111100;
DRAM[13201] = 8'b11111100;
DRAM[13202] = 8'b11111011;
DRAM[13203] = 8'b11111011;
DRAM[13204] = 8'b11111010;
DRAM[13205] = 8'b11111010;
DRAM[13206] = 8'b11111010;
DRAM[13207] = 8'b11111010;
DRAM[13208] = 8'b11111010;
DRAM[13209] = 8'b11111010;
DRAM[13210] = 8'b11111011;
DRAM[13211] = 8'b11111011;
DRAM[13212] = 8'b11111100;
DRAM[13213] = 8'b11111101;
DRAM[13214] = 8'b11111101;
DRAM[13215] = 8'b11111110;
DRAM[13216] = 8'b11111110;
DRAM[13217] = 8'b11111110;
DRAM[13218] = 8'b11111110;
DRAM[13219] = 8'b11111110;
DRAM[13220] = 8'b11111110;
DRAM[13221] = 8'b11111110;
DRAM[13222] = 8'b11111110;
DRAM[13223] = 8'b11111110;
DRAM[13224] = 8'b11111110;
DRAM[13225] = 8'b11111110;
DRAM[13226] = 8'b11111110;
DRAM[13227] = 8'b11111110;
DRAM[13228] = 8'b11111110;
DRAM[13229] = 8'b11111110;
DRAM[13230] = 8'b11111110;
DRAM[13231] = 8'b11111110;
DRAM[13232] = 8'b11111100;
DRAM[13233] = 8'b11111011;
DRAM[13234] = 8'b11111010;
DRAM[13235] = 8'b11111001;
DRAM[13236] = 8'b11110111;
DRAM[13237] = 8'b11110111;
DRAM[13238] = 8'b11111001;
DRAM[13239] = 8'b11111010;
DRAM[13240] = 8'b11111001;
DRAM[13241] = 8'b11111100;
DRAM[13242] = 8'b11111111;
DRAM[13243] = 8'b11111111;
DRAM[13244] = 8'b11111101;
DRAM[13245] = 8'b11111100;
DRAM[13246] = 8'b11111101;
DRAM[13247] = 8'b11111111;
DRAM[13248] = 8'b11111110;
DRAM[13249] = 8'b11111110;
DRAM[13250] = 8'b11111110;
DRAM[13251] = 8'b11111110;
DRAM[13252] = 8'b11111110;
DRAM[13253] = 8'b11111110;
DRAM[13254] = 8'b11111110;
DRAM[13255] = 8'b11111110;
DRAM[13256] = 8'b11111000;
DRAM[13257] = 8'b11111111;
DRAM[13258] = 8'b11111111;
DRAM[13259] = 8'b11111110;
DRAM[13260] = 8'b11111010;
DRAM[13261] = 8'b11111100;
DRAM[13262] = 8'b11111111;
DRAM[13263] = 8'b11111111;
DRAM[13264] = 8'b11111101;
DRAM[13265] = 8'b11100110;
DRAM[13266] = 8'b11010110;
DRAM[13267] = 8'b11000000;
DRAM[13268] = 8'b10011010;
DRAM[13269] = 8'b1111110;
DRAM[13270] = 8'b1111000;
DRAM[13271] = 8'b1111000;
DRAM[13272] = 8'b1101011;
DRAM[13273] = 8'b1100010;
DRAM[13274] = 8'b1011100;
DRAM[13275] = 8'b1011100;
DRAM[13276] = 8'b1011100;
DRAM[13277] = 8'b1011010;
DRAM[13278] = 8'b1011001;
DRAM[13279] = 8'b1011011;
DRAM[13280] = 8'b1011000;
DRAM[13281] = 8'b1011000;
DRAM[13282] = 8'b1010111;
DRAM[13283] = 8'b1010111;
DRAM[13284] = 8'b1010111;
DRAM[13285] = 8'b1010110;
DRAM[13286] = 8'b1010110;
DRAM[13287] = 8'b1010110;
DRAM[13288] = 8'b1010101;
DRAM[13289] = 8'b1010101;
DRAM[13290] = 8'b1010100;
DRAM[13291] = 8'b1010100;
DRAM[13292] = 8'b1010011;
DRAM[13293] = 8'b1010011;
DRAM[13294] = 8'b1010011;
DRAM[13295] = 8'b1010011;
DRAM[13296] = 8'b1010011;
DRAM[13297] = 8'b1010011;
DRAM[13298] = 8'b1010010;
DRAM[13299] = 8'b1010010;
DRAM[13300] = 8'b1010010;
DRAM[13301] = 8'b1010001;
DRAM[13302] = 8'b1010001;
DRAM[13303] = 8'b1010001;
DRAM[13304] = 8'b1010001;
DRAM[13305] = 8'b1010001;
DRAM[13306] = 8'b1010001;
DRAM[13307] = 8'b1010001;
DRAM[13308] = 8'b1010001;
DRAM[13309] = 8'b1010001;
DRAM[13310] = 8'b1010001;
DRAM[13311] = 8'b1010001;
DRAM[13312] = 8'b1100011;
DRAM[13313] = 8'b1100011;
DRAM[13314] = 8'b1100100;
DRAM[13315] = 8'b1100101;
DRAM[13316] = 8'b1100101;
DRAM[13317] = 8'b1100110;
DRAM[13318] = 8'b1100111;
DRAM[13319] = 8'b1100111;
DRAM[13320] = 8'b1101001;
DRAM[13321] = 8'b1101000;
DRAM[13322] = 8'b1100111;
DRAM[13323] = 8'b1100110;
DRAM[13324] = 8'b1100110;
DRAM[13325] = 8'b1101000;
DRAM[13326] = 8'b1101010;
DRAM[13327] = 8'b1101011;
DRAM[13328] = 8'b1101100;
DRAM[13329] = 8'b1101100;
DRAM[13330] = 8'b1101100;
DRAM[13331] = 8'b1101100;
DRAM[13332] = 8'b1101100;
DRAM[13333] = 8'b1101100;
DRAM[13334] = 8'b1101100;
DRAM[13335] = 8'b1101100;
DRAM[13336] = 8'b1101101;
DRAM[13337] = 8'b1101110;
DRAM[13338] = 8'b1101111;
DRAM[13339] = 8'b1110000;
DRAM[13340] = 8'b1110000;
DRAM[13341] = 8'b1110000;
DRAM[13342] = 8'b1110000;
DRAM[13343] = 8'b1101111;
DRAM[13344] = 8'b1110010;
DRAM[13345] = 8'b1110010;
DRAM[13346] = 8'b1110011;
DRAM[13347] = 8'b1110100;
DRAM[13348] = 8'b1110100;
DRAM[13349] = 8'b1110101;
DRAM[13350] = 8'b1110110;
DRAM[13351] = 8'b1110110;
DRAM[13352] = 8'b1110110;
DRAM[13353] = 8'b1110110;
DRAM[13354] = 8'b1110111;
DRAM[13355] = 8'b1111000;
DRAM[13356] = 8'b1111001;
DRAM[13357] = 8'b1111001;
DRAM[13358] = 8'b1111010;
DRAM[13359] = 8'b1111010;
DRAM[13360] = 8'b1111001;
DRAM[13361] = 8'b1111010;
DRAM[13362] = 8'b1111001;
DRAM[13363] = 8'b1111010;
DRAM[13364] = 8'b10000001;
DRAM[13365] = 8'b10001010;
DRAM[13366] = 8'b10001111;
DRAM[13367] = 8'b10001110;
DRAM[13368] = 8'b10001000;
DRAM[13369] = 8'b10010110;
DRAM[13370] = 8'b10100101;
DRAM[13371] = 8'b10110010;
DRAM[13372] = 8'b11000101;
DRAM[13373] = 8'b11100010;
DRAM[13374] = 8'b11111101;
DRAM[13375] = 8'b11111111;
DRAM[13376] = 8'b11111010;
DRAM[13377] = 8'b11111011;
DRAM[13378] = 8'b11111011;
DRAM[13379] = 8'b11111010;
DRAM[13380] = 8'b11111011;
DRAM[13381] = 8'b11111110;
DRAM[13382] = 8'b11111110;
DRAM[13383] = 8'b11111011;
DRAM[13384] = 8'b11111110;
DRAM[13385] = 8'b11111110;
DRAM[13386] = 8'b11111110;
DRAM[13387] = 8'b11111110;
DRAM[13388] = 8'b11111110;
DRAM[13389] = 8'b11111110;
DRAM[13390] = 8'b11111110;
DRAM[13391] = 8'b11111110;
DRAM[13392] = 8'b11111110;
DRAM[13393] = 8'b11111110;
DRAM[13394] = 8'b11111110;
DRAM[13395] = 8'b11111110;
DRAM[13396] = 8'b11111110;
DRAM[13397] = 8'b11111110;
DRAM[13398] = 8'b11111110;
DRAM[13399] = 8'b11111110;
DRAM[13400] = 8'b11111110;
DRAM[13401] = 8'b11111110;
DRAM[13402] = 8'b11111110;
DRAM[13403] = 8'b11111110;
DRAM[13404] = 8'b11111110;
DRAM[13405] = 8'b11111110;
DRAM[13406] = 8'b11111110;
DRAM[13407] = 8'b11111110;
DRAM[13408] = 8'b11111101;
DRAM[13409] = 8'b11111110;
DRAM[13410] = 8'b11111110;
DRAM[13411] = 8'b11111110;
DRAM[13412] = 8'b11111110;
DRAM[13413] = 8'b11111101;
DRAM[13414] = 8'b11111100;
DRAM[13415] = 8'b11111011;
DRAM[13416] = 8'b11111010;
DRAM[13417] = 8'b11111011;
DRAM[13418] = 8'b11111100;
DRAM[13419] = 8'b11111100;
DRAM[13420] = 8'b11111101;
DRAM[13421] = 8'b11111100;
DRAM[13422] = 8'b11111100;
DRAM[13423] = 8'b11111011;
DRAM[13424] = 8'b11111001;
DRAM[13425] = 8'b11111010;
DRAM[13426] = 8'b11111011;
DRAM[13427] = 8'b11111100;
DRAM[13428] = 8'b11111101;
DRAM[13429] = 8'b11111101;
DRAM[13430] = 8'b11111100;
DRAM[13431] = 8'b11111100;
DRAM[13432] = 8'b11111011;
DRAM[13433] = 8'b11111011;
DRAM[13434] = 8'b11111100;
DRAM[13435] = 8'b11111100;
DRAM[13436] = 8'b11111100;
DRAM[13437] = 8'b11111101;
DRAM[13438] = 8'b11111101;
DRAM[13439] = 8'b11111101;
DRAM[13440] = 8'b11111110;
DRAM[13441] = 8'b11111111;
DRAM[13442] = 8'b11111111;
DRAM[13443] = 8'b11111111;
DRAM[13444] = 8'b11111111;
DRAM[13445] = 8'b11111111;
DRAM[13446] = 8'b11111111;
DRAM[13447] = 8'b11111111;
DRAM[13448] = 8'b11111110;
DRAM[13449] = 8'b11111111;
DRAM[13450] = 8'b11111111;
DRAM[13451] = 8'b11111111;
DRAM[13452] = 8'b11111110;
DRAM[13453] = 8'b11111110;
DRAM[13454] = 8'b11111100;
DRAM[13455] = 8'b11111100;
DRAM[13456] = 8'b11111011;
DRAM[13457] = 8'b11111011;
DRAM[13458] = 8'b11111001;
DRAM[13459] = 8'b11111000;
DRAM[13460] = 8'b11111000;
DRAM[13461] = 8'b11111000;
DRAM[13462] = 8'b11111001;
DRAM[13463] = 8'b11111001;
DRAM[13464] = 8'b11111000;
DRAM[13465] = 8'b11111001;
DRAM[13466] = 8'b11111001;
DRAM[13467] = 8'b11111010;
DRAM[13468] = 8'b11111011;
DRAM[13469] = 8'b11111100;
DRAM[13470] = 8'b11111101;
DRAM[13471] = 8'b11111101;
DRAM[13472] = 8'b11111110;
DRAM[13473] = 8'b11111110;
DRAM[13474] = 8'b11111110;
DRAM[13475] = 8'b11111110;
DRAM[13476] = 8'b11111110;
DRAM[13477] = 8'b11111110;
DRAM[13478] = 8'b11111110;
DRAM[13479] = 8'b11111110;
DRAM[13480] = 8'b11111100;
DRAM[13481] = 8'b11111100;
DRAM[13482] = 8'b11111100;
DRAM[13483] = 8'b11111100;
DRAM[13484] = 8'b11111100;
DRAM[13485] = 8'b11111100;
DRAM[13486] = 8'b11111100;
DRAM[13487] = 8'b11111100;
DRAM[13488] = 8'b11111001;
DRAM[13489] = 8'b11111100;
DRAM[13490] = 8'b11111110;
DRAM[13491] = 8'b11111010;
DRAM[13492] = 8'b11110010;
DRAM[13493] = 8'b11101110;
DRAM[13494] = 8'b11110000;
DRAM[13495] = 8'b11110101;
DRAM[13496] = 8'b11111000;
DRAM[13497] = 8'b11111011;
DRAM[13498] = 8'b11111110;
DRAM[13499] = 8'b11111111;
DRAM[13500] = 8'b11111111;
DRAM[13501] = 8'b11111110;
DRAM[13502] = 8'b11111100;
DRAM[13503] = 8'b11111010;
DRAM[13504] = 8'b11111110;
DRAM[13505] = 8'b11111110;
DRAM[13506] = 8'b11111110;
DRAM[13507] = 8'b11111110;
DRAM[13508] = 8'b11111110;
DRAM[13509] = 8'b11111110;
DRAM[13510] = 8'b11111110;
DRAM[13511] = 8'b11111110;
DRAM[13512] = 8'b11111011;
DRAM[13513] = 8'b11111111;
DRAM[13514] = 8'b11111111;
DRAM[13515] = 8'b11111110;
DRAM[13516] = 8'b11111011;
DRAM[13517] = 8'b11111010;
DRAM[13518] = 8'b11111000;
DRAM[13519] = 8'b11110110;
DRAM[13520] = 8'b11111011;
DRAM[13521] = 8'b11110010;
DRAM[13522] = 8'b11110000;
DRAM[13523] = 8'b11011111;
DRAM[13524] = 8'b10110101;
DRAM[13525] = 8'b10010001;
DRAM[13526] = 8'b10000001;
DRAM[13527] = 8'b1111011;
DRAM[13528] = 8'b1110110;
DRAM[13529] = 8'b1101010;
DRAM[13530] = 8'b1100000;
DRAM[13531] = 8'b1011101;
DRAM[13532] = 8'b1011110;
DRAM[13533] = 8'b1011101;
DRAM[13534] = 8'b1011101;
DRAM[13535] = 8'b1011111;
DRAM[13536] = 8'b1011000;
DRAM[13537] = 8'b1011000;
DRAM[13538] = 8'b1011000;
DRAM[13539] = 8'b1010111;
DRAM[13540] = 8'b1010111;
DRAM[13541] = 8'b1010111;
DRAM[13542] = 8'b1010110;
DRAM[13543] = 8'b1010110;
DRAM[13544] = 8'b1010101;
DRAM[13545] = 8'b1010101;
DRAM[13546] = 8'b1010101;
DRAM[13547] = 8'b1010100;
DRAM[13548] = 8'b1010100;
DRAM[13549] = 8'b1010100;
DRAM[13550] = 8'b1010011;
DRAM[13551] = 8'b1010011;
DRAM[13552] = 8'b1010011;
DRAM[13553] = 8'b1010011;
DRAM[13554] = 8'b1010011;
DRAM[13555] = 8'b1010010;
DRAM[13556] = 8'b1010010;
DRAM[13557] = 8'b1010010;
DRAM[13558] = 8'b1010001;
DRAM[13559] = 8'b1010001;
DRAM[13560] = 8'b1010001;
DRAM[13561] = 8'b1010001;
DRAM[13562] = 8'b1010001;
DRAM[13563] = 8'b1010001;
DRAM[13564] = 8'b1010001;
DRAM[13565] = 8'b1010001;
DRAM[13566] = 8'b1010001;
DRAM[13567] = 8'b1010001;
DRAM[13568] = 8'b1100011;
DRAM[13569] = 8'b1100011;
DRAM[13570] = 8'b1100100;
DRAM[13571] = 8'b1100101;
DRAM[13572] = 8'b1100101;
DRAM[13573] = 8'b1100110;
DRAM[13574] = 8'b1100111;
DRAM[13575] = 8'b1100111;
DRAM[13576] = 8'b1101000;
DRAM[13577] = 8'b1100111;
DRAM[13578] = 8'b1100111;
DRAM[13579] = 8'b1100111;
DRAM[13580] = 8'b1101000;
DRAM[13581] = 8'b1101000;
DRAM[13582] = 8'b1101001;
DRAM[13583] = 8'b1101010;
DRAM[13584] = 8'b1101011;
DRAM[13585] = 8'b1101011;
DRAM[13586] = 8'b1101011;
DRAM[13587] = 8'b1101100;
DRAM[13588] = 8'b1101100;
DRAM[13589] = 8'b1101101;
DRAM[13590] = 8'b1101101;
DRAM[13591] = 8'b1101101;
DRAM[13592] = 8'b1101101;
DRAM[13593] = 8'b1101110;
DRAM[13594] = 8'b1101111;
DRAM[13595] = 8'b1110000;
DRAM[13596] = 8'b1110000;
DRAM[13597] = 8'b1110000;
DRAM[13598] = 8'b1110000;
DRAM[13599] = 8'b1101111;
DRAM[13600] = 8'b1110010;
DRAM[13601] = 8'b1110010;
DRAM[13602] = 8'b1110011;
DRAM[13603] = 8'b1110100;
DRAM[13604] = 8'b1110100;
DRAM[13605] = 8'b1110101;
DRAM[13606] = 8'b1110110;
DRAM[13607] = 8'b1110110;
DRAM[13608] = 8'b1110111;
DRAM[13609] = 8'b1110111;
DRAM[13610] = 8'b1110111;
DRAM[13611] = 8'b1111000;
DRAM[13612] = 8'b1111001;
DRAM[13613] = 8'b1111010;
DRAM[13614] = 8'b1111010;
DRAM[13615] = 8'b1111011;
DRAM[13616] = 8'b1111100;
DRAM[13617] = 8'b1111100;
DRAM[13618] = 8'b1111110;
DRAM[13619] = 8'b10000001;
DRAM[13620] = 8'b10000001;
DRAM[13621] = 8'b10000000;
DRAM[13622] = 8'b10000101;
DRAM[13623] = 8'b10001100;
DRAM[13624] = 8'b10001010;
DRAM[13625] = 8'b10101100;
DRAM[13626] = 8'b11010100;
DRAM[13627] = 8'b11101100;
DRAM[13628] = 8'b11111001;
DRAM[13629] = 8'b11111101;
DRAM[13630] = 8'b11111001;
DRAM[13631] = 8'b11110000;
DRAM[13632] = 8'b11111101;
DRAM[13633] = 8'b11111100;
DRAM[13634] = 8'b11111010;
DRAM[13635] = 8'b11111010;
DRAM[13636] = 8'b11111011;
DRAM[13637] = 8'b11111101;
DRAM[13638] = 8'b11111101;
DRAM[13639] = 8'b11111100;
DRAM[13640] = 8'b11111111;
DRAM[13641] = 8'b11111111;
DRAM[13642] = 8'b11111110;
DRAM[13643] = 8'b11111110;
DRAM[13644] = 8'b11111110;
DRAM[13645] = 8'b11111110;
DRAM[13646] = 8'b11111101;
DRAM[13647] = 8'b11111101;
DRAM[13648] = 8'b11111101;
DRAM[13649] = 8'b11111101;
DRAM[13650] = 8'b11111101;
DRAM[13651] = 8'b11111101;
DRAM[13652] = 8'b11111101;
DRAM[13653] = 8'b11111101;
DRAM[13654] = 8'b11111101;
DRAM[13655] = 8'b11111101;
DRAM[13656] = 8'b11111101;
DRAM[13657] = 8'b11111101;
DRAM[13658] = 8'b11111101;
DRAM[13659] = 8'b11111101;
DRAM[13660] = 8'b11111101;
DRAM[13661] = 8'b11111101;
DRAM[13662] = 8'b11111101;
DRAM[13663] = 8'b11111101;
DRAM[13664] = 8'b11111101;
DRAM[13665] = 8'b11111110;
DRAM[13666] = 8'b11111110;
DRAM[13667] = 8'b11111110;
DRAM[13668] = 8'b11111110;
DRAM[13669] = 8'b11111101;
DRAM[13670] = 8'b11111100;
DRAM[13671] = 8'b11111011;
DRAM[13672] = 8'b11111010;
DRAM[13673] = 8'b11111011;
DRAM[13674] = 8'b11111011;
DRAM[13675] = 8'b11111100;
DRAM[13676] = 8'b11111100;
DRAM[13677] = 8'b11111011;
DRAM[13678] = 8'b11111010;
DRAM[13679] = 8'b11111010;
DRAM[13680] = 8'b11110111;
DRAM[13681] = 8'b11111001;
DRAM[13682] = 8'b11111010;
DRAM[13683] = 8'b11111100;
DRAM[13684] = 8'b11111101;
DRAM[13685] = 8'b11111101;
DRAM[13686] = 8'b11111100;
DRAM[13687] = 8'b11111011;
DRAM[13688] = 8'b11111011;
DRAM[13689] = 8'b11111011;
DRAM[13690] = 8'b11111011;
DRAM[13691] = 8'b11111100;
DRAM[13692] = 8'b11111100;
DRAM[13693] = 8'b11111101;
DRAM[13694] = 8'b11111101;
DRAM[13695] = 8'b11111101;
DRAM[13696] = 8'b11111101;
DRAM[13697] = 8'b11111110;
DRAM[13698] = 8'b11111111;
DRAM[13699] = 8'b11111111;
DRAM[13700] = 8'b11111111;
DRAM[13701] = 8'b11111111;
DRAM[13702] = 8'b11111111;
DRAM[13703] = 8'b11111111;
DRAM[13704] = 8'b11111110;
DRAM[13705] = 8'b11111110;
DRAM[13706] = 8'b11111110;
DRAM[13707] = 8'b11111110;
DRAM[13708] = 8'b11111101;
DRAM[13709] = 8'b11111100;
DRAM[13710] = 8'b11111011;
DRAM[13711] = 8'b11111010;
DRAM[13712] = 8'b11111010;
DRAM[13713] = 8'b11111001;
DRAM[13714] = 8'b11110111;
DRAM[13715] = 8'b11110110;
DRAM[13716] = 8'b11110101;
DRAM[13717] = 8'b11110110;
DRAM[13718] = 8'b11110111;
DRAM[13719] = 8'b11111000;
DRAM[13720] = 8'b11110110;
DRAM[13721] = 8'b11110110;
DRAM[13722] = 8'b11110111;
DRAM[13723] = 8'b11111000;
DRAM[13724] = 8'b11111001;
DRAM[13725] = 8'b11111010;
DRAM[13726] = 8'b11111011;
DRAM[13727] = 8'b11111100;
DRAM[13728] = 8'b11111101;
DRAM[13729] = 8'b11111101;
DRAM[13730] = 8'b11111101;
DRAM[13731] = 8'b11111101;
DRAM[13732] = 8'b11111101;
DRAM[13733] = 8'b11111101;
DRAM[13734] = 8'b11111101;
DRAM[13735] = 8'b11111101;
DRAM[13736] = 8'b11111100;
DRAM[13737] = 8'b11111100;
DRAM[13738] = 8'b11111100;
DRAM[13739] = 8'b11111011;
DRAM[13740] = 8'b11111011;
DRAM[13741] = 8'b11111011;
DRAM[13742] = 8'b11111010;
DRAM[13743] = 8'b11111010;
DRAM[13744] = 8'b11111001;
DRAM[13745] = 8'b11111110;
DRAM[13746] = 8'b11111111;
DRAM[13747] = 8'b11111100;
DRAM[13748] = 8'b11110010;
DRAM[13749] = 8'b11101011;
DRAM[13750] = 8'b11101011;
DRAM[13751] = 8'b11101101;
DRAM[13752] = 8'b11110000;
DRAM[13753] = 8'b11110001;
DRAM[13754] = 8'b11110100;
DRAM[13755] = 8'b11111010;
DRAM[13756] = 8'b11111111;
DRAM[13757] = 8'b11111111;
DRAM[13758] = 8'b11111101;
DRAM[13759] = 8'b11111001;
DRAM[13760] = 8'b11111110;
DRAM[13761] = 8'b11111110;
DRAM[13762] = 8'b11111110;
DRAM[13763] = 8'b11111110;
DRAM[13764] = 8'b11111110;
DRAM[13765] = 8'b11111110;
DRAM[13766] = 8'b11111110;
DRAM[13767] = 8'b11111110;
DRAM[13768] = 8'b11111111;
DRAM[13769] = 8'b11111111;
DRAM[13770] = 8'b11111100;
DRAM[13771] = 8'b11111010;
DRAM[13772] = 8'b11111010;
DRAM[13773] = 8'b11111011;
DRAM[13774] = 8'b11111010;
DRAM[13775] = 8'b11111000;
DRAM[13776] = 8'b11111111;
DRAM[13777] = 8'b11111011;
DRAM[13778] = 8'b11111001;
DRAM[13779] = 8'b11110011;
DRAM[13780] = 8'b11011110;
DRAM[13781] = 8'b11001010;
DRAM[13782] = 8'b10110101;
DRAM[13783] = 8'b10011111;
DRAM[13784] = 8'b10000111;
DRAM[13785] = 8'b1111001;
DRAM[13786] = 8'b1101100;
DRAM[13787] = 8'b1100111;
DRAM[13788] = 8'b1100101;
DRAM[13789] = 8'b1100010;
DRAM[13790] = 8'b1100000;
DRAM[13791] = 8'b1100000;
DRAM[13792] = 8'b1011001;
DRAM[13793] = 8'b1011000;
DRAM[13794] = 8'b1011000;
DRAM[13795] = 8'b1011000;
DRAM[13796] = 8'b1010111;
DRAM[13797] = 8'b1010111;
DRAM[13798] = 8'b1010111;
DRAM[13799] = 8'b1010111;
DRAM[13800] = 8'b1011000;
DRAM[13801] = 8'b1011000;
DRAM[13802] = 8'b1010111;
DRAM[13803] = 8'b1010111;
DRAM[13804] = 8'b1010111;
DRAM[13805] = 8'b1010110;
DRAM[13806] = 8'b1010110;
DRAM[13807] = 8'b1010110;
DRAM[13808] = 8'b1010100;
DRAM[13809] = 8'b1010011;
DRAM[13810] = 8'b1010011;
DRAM[13811] = 8'b1010011;
DRAM[13812] = 8'b1010010;
DRAM[13813] = 8'b1010010;
DRAM[13814] = 8'b1010010;
DRAM[13815] = 8'b1010010;
DRAM[13816] = 8'b1010010;
DRAM[13817] = 8'b1010010;
DRAM[13818] = 8'b1010010;
DRAM[13819] = 8'b1010010;
DRAM[13820] = 8'b1010010;
DRAM[13821] = 8'b1010010;
DRAM[13822] = 8'b1010010;
DRAM[13823] = 8'b1010010;
DRAM[13824] = 8'b1100011;
DRAM[13825] = 8'b1100011;
DRAM[13826] = 8'b1100100;
DRAM[13827] = 8'b1100101;
DRAM[13828] = 8'b1100101;
DRAM[13829] = 8'b1100110;
DRAM[13830] = 8'b1100111;
DRAM[13831] = 8'b1100111;
DRAM[13832] = 8'b1100110;
DRAM[13833] = 8'b1100111;
DRAM[13834] = 8'b1101000;
DRAM[13835] = 8'b1101000;
DRAM[13836] = 8'b1101001;
DRAM[13837] = 8'b1101001;
DRAM[13838] = 8'b1101001;
DRAM[13839] = 8'b1101000;
DRAM[13840] = 8'b1101001;
DRAM[13841] = 8'b1101010;
DRAM[13842] = 8'b1101010;
DRAM[13843] = 8'b1101011;
DRAM[13844] = 8'b1101101;
DRAM[13845] = 8'b1101110;
DRAM[13846] = 8'b1101110;
DRAM[13847] = 8'b1101111;
DRAM[13848] = 8'b1101101;
DRAM[13849] = 8'b1101110;
DRAM[13850] = 8'b1101111;
DRAM[13851] = 8'b1110000;
DRAM[13852] = 8'b1110000;
DRAM[13853] = 8'b1110000;
DRAM[13854] = 8'b1110000;
DRAM[13855] = 8'b1101111;
DRAM[13856] = 8'b1110010;
DRAM[13857] = 8'b1110010;
DRAM[13858] = 8'b1110011;
DRAM[13859] = 8'b1110100;
DRAM[13860] = 8'b1110100;
DRAM[13861] = 8'b1110101;
DRAM[13862] = 8'b1110110;
DRAM[13863] = 8'b1110110;
DRAM[13864] = 8'b1110111;
DRAM[13865] = 8'b1110111;
DRAM[13866] = 8'b1111000;
DRAM[13867] = 8'b1111000;
DRAM[13868] = 8'b1111001;
DRAM[13869] = 8'b1111010;
DRAM[13870] = 8'b1111011;
DRAM[13871] = 8'b1111011;
DRAM[13872] = 8'b1111110;
DRAM[13873] = 8'b1111101;
DRAM[13874] = 8'b10000001;
DRAM[13875] = 8'b10000100;
DRAM[13876] = 8'b1111011;
DRAM[13877] = 8'b1110110;
DRAM[13878] = 8'b10001011;
DRAM[13879] = 8'b10101000;
DRAM[13880] = 8'b11011010;
DRAM[13881] = 8'b11101110;
DRAM[13882] = 8'b11111100;
DRAM[13883] = 8'b11111100;
DRAM[13884] = 8'b11111001;
DRAM[13885] = 8'b11111101;
DRAM[13886] = 8'b11111111;
DRAM[13887] = 8'b11111100;
DRAM[13888] = 8'b11111110;
DRAM[13889] = 8'b11111101;
DRAM[13890] = 8'b11111100;
DRAM[13891] = 8'b11111101;
DRAM[13892] = 8'b11111101;
DRAM[13893] = 8'b11111101;
DRAM[13894] = 8'b11111101;
DRAM[13895] = 8'b11111110;
DRAM[13896] = 8'b11111111;
DRAM[13897] = 8'b11111111;
DRAM[13898] = 8'b11111111;
DRAM[13899] = 8'b11111110;
DRAM[13900] = 8'b11111110;
DRAM[13901] = 8'b11111101;
DRAM[13902] = 8'b11111101;
DRAM[13903] = 8'b11111101;
DRAM[13904] = 8'b11111101;
DRAM[13905] = 8'b11111101;
DRAM[13906] = 8'b11111101;
DRAM[13907] = 8'b11111101;
DRAM[13908] = 8'b11111101;
DRAM[13909] = 8'b11111101;
DRAM[13910] = 8'b11111101;
DRAM[13911] = 8'b11111101;
DRAM[13912] = 8'b11111101;
DRAM[13913] = 8'b11111101;
DRAM[13914] = 8'b11111101;
DRAM[13915] = 8'b11111101;
DRAM[13916] = 8'b11111101;
DRAM[13917] = 8'b11111101;
DRAM[13918] = 8'b11111101;
DRAM[13919] = 8'b11111101;
DRAM[13920] = 8'b11111101;
DRAM[13921] = 8'b11111110;
DRAM[13922] = 8'b11111110;
DRAM[13923] = 8'b11111110;
DRAM[13924] = 8'b11111110;
DRAM[13925] = 8'b11111101;
DRAM[13926] = 8'b11111100;
DRAM[13927] = 8'b11111011;
DRAM[13928] = 8'b11111011;
DRAM[13929] = 8'b11111011;
DRAM[13930] = 8'b11111100;
DRAM[13931] = 8'b11111011;
DRAM[13932] = 8'b11111011;
DRAM[13933] = 8'b11111010;
DRAM[13934] = 8'b11111000;
DRAM[13935] = 8'b11111000;
DRAM[13936] = 8'b11110110;
DRAM[13937] = 8'b11110111;
DRAM[13938] = 8'b11111010;
DRAM[13939] = 8'b11111100;
DRAM[13940] = 8'b11111101;
DRAM[13941] = 8'b11111100;
DRAM[13942] = 8'b11111011;
DRAM[13943] = 8'b11111010;
DRAM[13944] = 8'b11111001;
DRAM[13945] = 8'b11111010;
DRAM[13946] = 8'b11111010;
DRAM[13947] = 8'b11111010;
DRAM[13948] = 8'b11111011;
DRAM[13949] = 8'b11111011;
DRAM[13950] = 8'b11111011;
DRAM[13951] = 8'b11111100;
DRAM[13952] = 8'b11111010;
DRAM[13953] = 8'b11111011;
DRAM[13954] = 8'b11111101;
DRAM[13955] = 8'b11111110;
DRAM[13956] = 8'b11111110;
DRAM[13957] = 8'b11111110;
DRAM[13958] = 8'b11111101;
DRAM[13959] = 8'b11111101;
DRAM[13960] = 8'b11111101;
DRAM[13961] = 8'b11111101;
DRAM[13962] = 8'b11111101;
DRAM[13963] = 8'b11111101;
DRAM[13964] = 8'b11111100;
DRAM[13965] = 8'b11111011;
DRAM[13966] = 8'b11111001;
DRAM[13967] = 8'b11111001;
DRAM[13968] = 8'b11111000;
DRAM[13969] = 8'b11110111;
DRAM[13970] = 8'b11110101;
DRAM[13971] = 8'b11110011;
DRAM[13972] = 8'b11110011;
DRAM[13973] = 8'b11110100;
DRAM[13974] = 8'b11110101;
DRAM[13975] = 8'b11110110;
DRAM[13976] = 8'b11110100;
DRAM[13977] = 8'b11110100;
DRAM[13978] = 8'b11110101;
DRAM[13979] = 8'b11110110;
DRAM[13980] = 8'b11111000;
DRAM[13981] = 8'b11111001;
DRAM[13982] = 8'b11111010;
DRAM[13983] = 8'b11111010;
DRAM[13984] = 8'b11111101;
DRAM[13985] = 8'b11111101;
DRAM[13986] = 8'b11111101;
DRAM[13987] = 8'b11111101;
DRAM[13988] = 8'b11111101;
DRAM[13989] = 8'b11111101;
DRAM[13990] = 8'b11111101;
DRAM[13991] = 8'b11111101;
DRAM[13992] = 8'b11111101;
DRAM[13993] = 8'b11111101;
DRAM[13994] = 8'b11111101;
DRAM[13995] = 8'b11111100;
DRAM[13996] = 8'b11111100;
DRAM[13997] = 8'b11111011;
DRAM[13998] = 8'b11111011;
DRAM[13999] = 8'b11111011;
DRAM[14000] = 8'b11111101;
DRAM[14001] = 8'b11111101;
DRAM[14002] = 8'b11111101;
DRAM[14003] = 8'b11111100;
DRAM[14004] = 8'b11111000;
DRAM[14005] = 8'b11110010;
DRAM[14006] = 8'b11101011;
DRAM[14007] = 8'b11100110;
DRAM[14008] = 8'b11011111;
DRAM[14009] = 8'b11011100;
DRAM[14010] = 8'b11011100;
DRAM[14011] = 8'b11100110;
DRAM[14012] = 8'b11110101;
DRAM[14013] = 8'b11111111;
DRAM[14014] = 8'b11111110;
DRAM[14015] = 8'b11111010;
DRAM[14016] = 8'b11111110;
DRAM[14017] = 8'b11111110;
DRAM[14018] = 8'b11111110;
DRAM[14019] = 8'b11111110;
DRAM[14020] = 8'b11111110;
DRAM[14021] = 8'b11111110;
DRAM[14022] = 8'b11111110;
DRAM[14023] = 8'b11111110;
DRAM[14024] = 8'b11111111;
DRAM[14025] = 8'b11111111;
DRAM[14026] = 8'b11111011;
DRAM[14027] = 8'b11111011;
DRAM[14028] = 8'b11111100;
DRAM[14029] = 8'b11111101;
DRAM[14030] = 8'b11111110;
DRAM[14031] = 8'b11111110;
DRAM[14032] = 8'b11111001;
DRAM[14033] = 8'b11110100;
DRAM[14034] = 8'b11110101;
DRAM[14035] = 8'b11110100;
DRAM[14036] = 8'b11110010;
DRAM[14037] = 8'b11110010;
DRAM[14038] = 8'b11100010;
DRAM[14039] = 8'b11000100;
DRAM[14040] = 8'b10011001;
DRAM[14041] = 8'b10001011;
DRAM[14042] = 8'b1111110;
DRAM[14043] = 8'b1110111;
DRAM[14044] = 8'b1110010;
DRAM[14045] = 8'b1101001;
DRAM[14046] = 8'b1100000;
DRAM[14047] = 8'b1011100;
DRAM[14048] = 8'b1011001;
DRAM[14049] = 8'b1011001;
DRAM[14050] = 8'b1011000;
DRAM[14051] = 8'b1011000;
DRAM[14052] = 8'b1011000;
DRAM[14053] = 8'b1010111;
DRAM[14054] = 8'b1010111;
DRAM[14055] = 8'b1010111;
DRAM[14056] = 8'b1011000;
DRAM[14057] = 8'b1011000;
DRAM[14058] = 8'b1011000;
DRAM[14059] = 8'b1010111;
DRAM[14060] = 8'b1010111;
DRAM[14061] = 8'b1010110;
DRAM[14062] = 8'b1010110;
DRAM[14063] = 8'b1010110;
DRAM[14064] = 8'b1010100;
DRAM[14065] = 8'b1010100;
DRAM[14066] = 8'b1010011;
DRAM[14067] = 8'b1010011;
DRAM[14068] = 8'b1010011;
DRAM[14069] = 8'b1010010;
DRAM[14070] = 8'b1010010;
DRAM[14071] = 8'b1010010;
DRAM[14072] = 8'b1010010;
DRAM[14073] = 8'b1010010;
DRAM[14074] = 8'b1010010;
DRAM[14075] = 8'b1010010;
DRAM[14076] = 8'b1010010;
DRAM[14077] = 8'b1010010;
DRAM[14078] = 8'b1010010;
DRAM[14079] = 8'b1010010;
DRAM[14080] = 8'b1100011;
DRAM[14081] = 8'b1100011;
DRAM[14082] = 8'b1100100;
DRAM[14083] = 8'b1100101;
DRAM[14084] = 8'b1100101;
DRAM[14085] = 8'b1100110;
DRAM[14086] = 8'b1100111;
DRAM[14087] = 8'b1100111;
DRAM[14088] = 8'b1100101;
DRAM[14089] = 8'b1100110;
DRAM[14090] = 8'b1101000;
DRAM[14091] = 8'b1101010;
DRAM[14092] = 8'b1101010;
DRAM[14093] = 8'b1101001;
DRAM[14094] = 8'b1101000;
DRAM[14095] = 8'b1100111;
DRAM[14096] = 8'b1101000;
DRAM[14097] = 8'b1101001;
DRAM[14098] = 8'b1101010;
DRAM[14099] = 8'b1101011;
DRAM[14100] = 8'b1101101;
DRAM[14101] = 8'b1101110;
DRAM[14102] = 8'b1101111;
DRAM[14103] = 8'b1110000;
DRAM[14104] = 8'b1101101;
DRAM[14105] = 8'b1101110;
DRAM[14106] = 8'b1101111;
DRAM[14107] = 8'b1110000;
DRAM[14108] = 8'b1110000;
DRAM[14109] = 8'b1110000;
DRAM[14110] = 8'b1110000;
DRAM[14111] = 8'b1101111;
DRAM[14112] = 8'b1110010;
DRAM[14113] = 8'b1110010;
DRAM[14114] = 8'b1110011;
DRAM[14115] = 8'b1110100;
DRAM[14116] = 8'b1110100;
DRAM[14117] = 8'b1110101;
DRAM[14118] = 8'b1110110;
DRAM[14119] = 8'b1110110;
DRAM[14120] = 8'b1110111;
DRAM[14121] = 8'b1110111;
DRAM[14122] = 8'b1111000;
DRAM[14123] = 8'b1111001;
DRAM[14124] = 8'b1111001;
DRAM[14125] = 8'b1111010;
DRAM[14126] = 8'b1111011;
DRAM[14127] = 8'b1111011;
DRAM[14128] = 8'b1111010;
DRAM[14129] = 8'b1111000;
DRAM[14130] = 8'b1111111;
DRAM[14131] = 8'b10000011;
DRAM[14132] = 8'b1111010;
DRAM[14133] = 8'b1111110;
DRAM[14134] = 8'b10101011;
DRAM[14135] = 8'b11100000;
DRAM[14136] = 8'b11101010;
DRAM[14137] = 8'b11111001;
DRAM[14138] = 8'b11111111;
DRAM[14139] = 8'b11111000;
DRAM[14140] = 8'b11110011;
DRAM[14141] = 8'b11111010;
DRAM[14142] = 8'b11111111;
DRAM[14143] = 8'b11111111;
DRAM[14144] = 8'b11111111;
DRAM[14145] = 8'b11111111;
DRAM[14146] = 8'b11111111;
DRAM[14147] = 8'b11111111;
DRAM[14148] = 8'b11111111;
DRAM[14149] = 8'b11111101;
DRAM[14150] = 8'b11111101;
DRAM[14151] = 8'b11111111;
DRAM[14152] = 8'b11111111;
DRAM[14153] = 8'b11111111;
DRAM[14154] = 8'b11111111;
DRAM[14155] = 8'b11111110;
DRAM[14156] = 8'b11111110;
DRAM[14157] = 8'b11111101;
DRAM[14158] = 8'b11111101;
DRAM[14159] = 8'b11111101;
DRAM[14160] = 8'b11111101;
DRAM[14161] = 8'b11111101;
DRAM[14162] = 8'b11111101;
DRAM[14163] = 8'b11111101;
DRAM[14164] = 8'b11111101;
DRAM[14165] = 8'b11111101;
DRAM[14166] = 8'b11111101;
DRAM[14167] = 8'b11111101;
DRAM[14168] = 8'b11111101;
DRAM[14169] = 8'b11111101;
DRAM[14170] = 8'b11111101;
DRAM[14171] = 8'b11111101;
DRAM[14172] = 8'b11111101;
DRAM[14173] = 8'b11111101;
DRAM[14174] = 8'b11111101;
DRAM[14175] = 8'b11111101;
DRAM[14176] = 8'b11111101;
DRAM[14177] = 8'b11111110;
DRAM[14178] = 8'b11111110;
DRAM[14179] = 8'b11111110;
DRAM[14180] = 8'b11111110;
DRAM[14181] = 8'b11111101;
DRAM[14182] = 8'b11111100;
DRAM[14183] = 8'b11111011;
DRAM[14184] = 8'b11111100;
DRAM[14185] = 8'b11111100;
DRAM[14186] = 8'b11111100;
DRAM[14187] = 8'b11111011;
DRAM[14188] = 8'b11111010;
DRAM[14189] = 8'b11111001;
DRAM[14190] = 8'b11110111;
DRAM[14191] = 8'b11110110;
DRAM[14192] = 8'b11110101;
DRAM[14193] = 8'b11110111;
DRAM[14194] = 8'b11111010;
DRAM[14195] = 8'b11111100;
DRAM[14196] = 8'b11111101;
DRAM[14197] = 8'b11111100;
DRAM[14198] = 8'b11111011;
DRAM[14199] = 8'b11111010;
DRAM[14200] = 8'b11111000;
DRAM[14201] = 8'b11111000;
DRAM[14202] = 8'b11111000;
DRAM[14203] = 8'b11111001;
DRAM[14204] = 8'b11111001;
DRAM[14205] = 8'b11111001;
DRAM[14206] = 8'b11111010;
DRAM[14207] = 8'b11111010;
DRAM[14208] = 8'b11111000;
DRAM[14209] = 8'b11111001;
DRAM[14210] = 8'b11111011;
DRAM[14211] = 8'b11111100;
DRAM[14212] = 8'b11111101;
DRAM[14213] = 8'b11111100;
DRAM[14214] = 8'b11111011;
DRAM[14215] = 8'b11111010;
DRAM[14216] = 8'b11111100;
DRAM[14217] = 8'b11111101;
DRAM[14218] = 8'b11111101;
DRAM[14219] = 8'b11111100;
DRAM[14220] = 8'b11111011;
DRAM[14221] = 8'b11111010;
DRAM[14222] = 8'b11111000;
DRAM[14223] = 8'b11111000;
DRAM[14224] = 8'b11110111;
DRAM[14225] = 8'b11110110;
DRAM[14226] = 8'b11110011;
DRAM[14227] = 8'b11110001;
DRAM[14228] = 8'b11110001;
DRAM[14229] = 8'b11110010;
DRAM[14230] = 8'b11110100;
DRAM[14231] = 8'b11110101;
DRAM[14232] = 8'b11110010;
DRAM[14233] = 8'b11110011;
DRAM[14234] = 8'b11110100;
DRAM[14235] = 8'b11110101;
DRAM[14236] = 8'b11110110;
DRAM[14237] = 8'b11111000;
DRAM[14238] = 8'b11111001;
DRAM[14239] = 8'b11111001;
DRAM[14240] = 8'b11111101;
DRAM[14241] = 8'b11111101;
DRAM[14242] = 8'b11111101;
DRAM[14243] = 8'b11111101;
DRAM[14244] = 8'b11111101;
DRAM[14245] = 8'b11111101;
DRAM[14246] = 8'b11111101;
DRAM[14247] = 8'b11111101;
DRAM[14248] = 8'b11111110;
DRAM[14249] = 8'b11111110;
DRAM[14250] = 8'b11111110;
DRAM[14251] = 8'b11111101;
DRAM[14252] = 8'b11111101;
DRAM[14253] = 8'b11111100;
DRAM[14254] = 8'b11111100;
DRAM[14255] = 8'b11111100;
DRAM[14256] = 8'b11111111;
DRAM[14257] = 8'b11111101;
DRAM[14258] = 8'b11111010;
DRAM[14259] = 8'b11111100;
DRAM[14260] = 8'b11111110;
DRAM[14261] = 8'b11111001;
DRAM[14262] = 8'b11101101;
DRAM[14263] = 8'b11100010;
DRAM[14264] = 8'b11001111;
DRAM[14265] = 8'b11001001;
DRAM[14266] = 8'b11000111;
DRAM[14267] = 8'b11010100;
DRAM[14268] = 8'b11101001;
DRAM[14269] = 8'b11111010;
DRAM[14270] = 8'b11111101;
DRAM[14271] = 8'b11111010;
DRAM[14272] = 8'b11111110;
DRAM[14273] = 8'b11111110;
DRAM[14274] = 8'b11111110;
DRAM[14275] = 8'b11111110;
DRAM[14276] = 8'b11111110;
DRAM[14277] = 8'b11111110;
DRAM[14278] = 8'b11111110;
DRAM[14279] = 8'b11111110;
DRAM[14280] = 8'b11111110;
DRAM[14281] = 8'b11111101;
DRAM[14282] = 8'b11111101;
DRAM[14283] = 8'b11111111;
DRAM[14284] = 8'b11111111;
DRAM[14285] = 8'b11111111;
DRAM[14286] = 8'b11111110;
DRAM[14287] = 8'b11111111;
DRAM[14288] = 8'b11110111;
DRAM[14289] = 8'b11111100;
DRAM[14290] = 8'b11111111;
DRAM[14291] = 8'b11111110;
DRAM[14292] = 8'b11111010;
DRAM[14293] = 8'b11111111;
DRAM[14294] = 8'b11110110;
DRAM[14295] = 8'b11011001;
DRAM[14296] = 8'b10100101;
DRAM[14297] = 8'b10011000;
DRAM[14298] = 8'b10001011;
DRAM[14299] = 8'b10000011;
DRAM[14300] = 8'b1111100;
DRAM[14301] = 8'b1101110;
DRAM[14302] = 8'b1011111;
DRAM[14303] = 8'b1010111;
DRAM[14304] = 8'b1011001;
DRAM[14305] = 8'b1011001;
DRAM[14306] = 8'b1011001;
DRAM[14307] = 8'b1011000;
DRAM[14308] = 8'b1011000;
DRAM[14309] = 8'b1010111;
DRAM[14310] = 8'b1010111;
DRAM[14311] = 8'b1010111;
DRAM[14312] = 8'b1010110;
DRAM[14313] = 8'b1010110;
DRAM[14314] = 8'b1010101;
DRAM[14315] = 8'b1010101;
DRAM[14316] = 8'b1010101;
DRAM[14317] = 8'b1010100;
DRAM[14318] = 8'b1010100;
DRAM[14319] = 8'b1010100;
DRAM[14320] = 8'b1010100;
DRAM[14321] = 8'b1010100;
DRAM[14322] = 8'b1010100;
DRAM[14323] = 8'b1010011;
DRAM[14324] = 8'b1010011;
DRAM[14325] = 8'b1010010;
DRAM[14326] = 8'b1010010;
DRAM[14327] = 8'b1010010;
DRAM[14328] = 8'b1010010;
DRAM[14329] = 8'b1010010;
DRAM[14330] = 8'b1010010;
DRAM[14331] = 8'b1010010;
DRAM[14332] = 8'b1010010;
DRAM[14333] = 8'b1010010;
DRAM[14334] = 8'b1010010;
DRAM[14335] = 8'b1010010;
DRAM[14336] = 8'b1100011;
DRAM[14337] = 8'b1100011;
DRAM[14338] = 8'b1100100;
DRAM[14339] = 8'b1100100;
DRAM[14340] = 8'b1100100;
DRAM[14341] = 8'b1100100;
DRAM[14342] = 8'b1100101;
DRAM[14343] = 8'b1100101;
DRAM[14344] = 8'b1100100;
DRAM[14345] = 8'b1100101;
DRAM[14346] = 8'b1100110;
DRAM[14347] = 8'b1100111;
DRAM[14348] = 8'b1101001;
DRAM[14349] = 8'b1101010;
DRAM[14350] = 8'b1101011;
DRAM[14351] = 8'b1101011;
DRAM[14352] = 8'b1101010;
DRAM[14353] = 8'b1101010;
DRAM[14354] = 8'b1101011;
DRAM[14355] = 8'b1101100;
DRAM[14356] = 8'b1101100;
DRAM[14357] = 8'b1101101;
DRAM[14358] = 8'b1101110;
DRAM[14359] = 8'b1101110;
DRAM[14360] = 8'b1110000;
DRAM[14361] = 8'b1110000;
DRAM[14362] = 8'b1110000;
DRAM[14363] = 8'b1110001;
DRAM[14364] = 8'b1110001;
DRAM[14365] = 8'b1110010;
DRAM[14366] = 8'b1110010;
DRAM[14367] = 8'b1110010;
DRAM[14368] = 8'b1110010;
DRAM[14369] = 8'b1110010;
DRAM[14370] = 8'b1110011;
DRAM[14371] = 8'b1110100;
DRAM[14372] = 8'b1110100;
DRAM[14373] = 8'b1110101;
DRAM[14374] = 8'b1110110;
DRAM[14375] = 8'b1110110;
DRAM[14376] = 8'b1110110;
DRAM[14377] = 8'b1111110;
DRAM[14378] = 8'b1111010;
DRAM[14379] = 8'b1110011;
DRAM[14380] = 8'b1110110;
DRAM[14381] = 8'b1110100;
DRAM[14382] = 8'b1110011;
DRAM[14383] = 8'b1111010;
DRAM[14384] = 8'b1111110;
DRAM[14385] = 8'b1111011;
DRAM[14386] = 8'b1111101;
DRAM[14387] = 8'b10001000;
DRAM[14388] = 8'b10011010;
DRAM[14389] = 8'b10111001;
DRAM[14390] = 8'b11100100;
DRAM[14391] = 8'b11111111;
DRAM[14392] = 8'b11111100;
DRAM[14393] = 8'b11111100;
DRAM[14394] = 8'b11111100;
DRAM[14395] = 8'b11111101;
DRAM[14396] = 8'b11111101;
DRAM[14397] = 8'b11111110;
DRAM[14398] = 8'b11111110;
DRAM[14399] = 8'b11111110;
DRAM[14400] = 8'b11111111;
DRAM[14401] = 8'b11111111;
DRAM[14402] = 8'b11111111;
DRAM[14403] = 8'b11111111;
DRAM[14404] = 8'b11111111;
DRAM[14405] = 8'b11111111;
DRAM[14406] = 8'b11111111;
DRAM[14407] = 8'b11111111;
DRAM[14408] = 8'b11111110;
DRAM[14409] = 8'b11111100;
DRAM[14410] = 8'b11111100;
DRAM[14411] = 8'b11111111;
DRAM[14412] = 8'b11111111;
DRAM[14413] = 8'b11111111;
DRAM[14414] = 8'b11111110;
DRAM[14415] = 8'b11111101;
DRAM[14416] = 8'b11111011;
DRAM[14417] = 8'b11111011;
DRAM[14418] = 8'b11111010;
DRAM[14419] = 8'b11111000;
DRAM[14420] = 8'b11110111;
DRAM[14421] = 8'b11110110;
DRAM[14422] = 8'b11110011;
DRAM[14423] = 8'b11101110;
DRAM[14424] = 8'b11110000;
DRAM[14425] = 8'b11110110;
DRAM[14426] = 8'b11111000;
DRAM[14427] = 8'b11110101;
DRAM[14428] = 8'b11110101;
DRAM[14429] = 8'b11111001;
DRAM[14430] = 8'b11111100;
DRAM[14431] = 8'b11111100;
DRAM[14432] = 8'b11111101;
DRAM[14433] = 8'b11111111;
DRAM[14434] = 8'b11111111;
DRAM[14435] = 8'b11111001;
DRAM[14436] = 8'b11110110;
DRAM[14437] = 8'b11111010;
DRAM[14438] = 8'b11111110;
DRAM[14439] = 8'b11111111;
DRAM[14440] = 8'b11110110;
DRAM[14441] = 8'b11111100;
DRAM[14442] = 8'b11111111;
DRAM[14443] = 8'b11111010;
DRAM[14444] = 8'b11110110;
DRAM[14445] = 8'b11110101;
DRAM[14446] = 8'b11110011;
DRAM[14447] = 8'b11110001;
DRAM[14448] = 8'b11110000;
DRAM[14449] = 8'b11110110;
DRAM[14450] = 8'b11110110;
DRAM[14451] = 8'b11110011;
DRAM[14452] = 8'b11110110;
DRAM[14453] = 8'b11111101;
DRAM[14454] = 8'b11111100;
DRAM[14455] = 8'b11110101;
DRAM[14456] = 8'b11111000;
DRAM[14457] = 8'b11111110;
DRAM[14458] = 8'b11111111;
DRAM[14459] = 8'b11111010;
DRAM[14460] = 8'b11110110;
DRAM[14461] = 8'b11110110;
DRAM[14462] = 8'b11111000;
DRAM[14463] = 8'b11111000;
DRAM[14464] = 8'b11111001;
DRAM[14465] = 8'b11111010;
DRAM[14466] = 8'b11111010;
DRAM[14467] = 8'b11111010;
DRAM[14468] = 8'b11111001;
DRAM[14469] = 8'b11111000;
DRAM[14470] = 8'b11111001;
DRAM[14471] = 8'b11111010;
DRAM[14472] = 8'b11111000;
DRAM[14473] = 8'b11111011;
DRAM[14474] = 8'b11111100;
DRAM[14475] = 8'b11111011;
DRAM[14476] = 8'b11111100;
DRAM[14477] = 8'b11111010;
DRAM[14478] = 8'b11110010;
DRAM[14479] = 8'b11101001;
DRAM[14480] = 8'b11101011;
DRAM[14481] = 8'b11101101;
DRAM[14482] = 8'b11111001;
DRAM[14483] = 8'b11111010;
DRAM[14484] = 8'b11101101;
DRAM[14485] = 8'b11101101;
DRAM[14486] = 8'b11110110;
DRAM[14487] = 8'b11110111;
DRAM[14488] = 8'b11110110;
DRAM[14489] = 8'b11101111;
DRAM[14490] = 8'b11101110;
DRAM[14491] = 8'b11110110;
DRAM[14492] = 8'b11110111;
DRAM[14493] = 8'b11110001;
DRAM[14494] = 8'b11110011;
DRAM[14495] = 8'b11111101;
DRAM[14496] = 8'b11111010;
DRAM[14497] = 8'b11111000;
DRAM[14498] = 8'b11110111;
DRAM[14499] = 8'b11111001;
DRAM[14500] = 8'b11111101;
DRAM[14501] = 8'b11111111;
DRAM[14502] = 8'b11111111;
DRAM[14503] = 8'b11111100;
DRAM[14504] = 8'b11111011;
DRAM[14505] = 8'b11111111;
DRAM[14506] = 8'b11111111;
DRAM[14507] = 8'b11111101;
DRAM[14508] = 8'b11111001;
DRAM[14509] = 8'b11111101;
DRAM[14510] = 8'b11111111;
DRAM[14511] = 8'b11111111;
DRAM[14512] = 8'b11111000;
DRAM[14513] = 8'b11111110;
DRAM[14514] = 8'b11111101;
DRAM[14515] = 8'b11110110;
DRAM[14516] = 8'b11110111;
DRAM[14517] = 8'b11111100;
DRAM[14518] = 8'b11110111;
DRAM[14519] = 8'b11101011;
DRAM[14520] = 8'b11001010;
DRAM[14521] = 8'b11001011;
DRAM[14522] = 8'b11000111;
DRAM[14523] = 8'b11000011;
DRAM[14524] = 8'b11001111;
DRAM[14525] = 8'b11100111;
DRAM[14526] = 8'b11110111;
DRAM[14527] = 8'b11111001;
DRAM[14528] = 8'b11111111;
DRAM[14529] = 8'b11110100;
DRAM[14530] = 8'b11111101;
DRAM[14531] = 8'b11111111;
DRAM[14532] = 8'b11111001;
DRAM[14533] = 8'b11110110;
DRAM[14534] = 8'b11111111;
DRAM[14535] = 8'b11111101;
DRAM[14536] = 8'b11111110;
DRAM[14537] = 8'b11111111;
DRAM[14538] = 8'b11111111;
DRAM[14539] = 8'b11111111;
DRAM[14540] = 8'b11111101;
DRAM[14541] = 8'b11111100;
DRAM[14542] = 8'b11111101;
DRAM[14543] = 8'b11111110;
DRAM[14544] = 8'b11111011;
DRAM[14545] = 8'b11111001;
DRAM[14546] = 8'b11111001;
DRAM[14547] = 8'b11111010;
DRAM[14548] = 8'b11111100;
DRAM[14549] = 8'b11111011;
DRAM[14550] = 8'b11110110;
DRAM[14551] = 8'b11110010;
DRAM[14552] = 8'b11011101;
DRAM[14553] = 8'b10101101;
DRAM[14554] = 8'b10000011;
DRAM[14555] = 8'b1111010;
DRAM[14556] = 8'b1111010;
DRAM[14557] = 8'b1101111;
DRAM[14558] = 8'b1100100;
DRAM[14559] = 8'b1100011;
DRAM[14560] = 8'b1011101;
DRAM[14561] = 8'b1011101;
DRAM[14562] = 8'b1011011;
DRAM[14563] = 8'b1011000;
DRAM[14564] = 8'b1011000;
DRAM[14565] = 8'b1011010;
DRAM[14566] = 8'b1011001;
DRAM[14567] = 8'b1011000;
DRAM[14568] = 8'b1010110;
DRAM[14569] = 8'b1010111;
DRAM[14570] = 8'b1011000;
DRAM[14571] = 8'b1011001;
DRAM[14572] = 8'b1011000;
DRAM[14573] = 8'b1010111;
DRAM[14574] = 8'b1010101;
DRAM[14575] = 8'b1010100;
DRAM[14576] = 8'b1010011;
DRAM[14577] = 8'b1010100;
DRAM[14578] = 8'b1010101;
DRAM[14579] = 8'b1010110;
DRAM[14580] = 8'b1010101;
DRAM[14581] = 8'b1010100;
DRAM[14582] = 8'b1010010;
DRAM[14583] = 8'b1010001;
DRAM[14584] = 8'b1010101;
DRAM[14585] = 8'b1010100;
DRAM[14586] = 8'b1010011;
DRAM[14587] = 8'b1010010;
DRAM[14588] = 8'b1010010;
DRAM[14589] = 8'b1010010;
DRAM[14590] = 8'b1010010;
DRAM[14591] = 8'b1010011;
DRAM[14592] = 8'b1100011;
DRAM[14593] = 8'b1100011;
DRAM[14594] = 8'b1100100;
DRAM[14595] = 8'b1100100;
DRAM[14596] = 8'b1100100;
DRAM[14597] = 8'b1100101;
DRAM[14598] = 8'b1100101;
DRAM[14599] = 8'b1100101;
DRAM[14600] = 8'b1100101;
DRAM[14601] = 8'b1100101;
DRAM[14602] = 8'b1100110;
DRAM[14603] = 8'b1100111;
DRAM[14604] = 8'b1101001;
DRAM[14605] = 8'b1101010;
DRAM[14606] = 8'b1101011;
DRAM[14607] = 8'b1101011;
DRAM[14608] = 8'b1101010;
DRAM[14609] = 8'b1101010;
DRAM[14610] = 8'b1101011;
DRAM[14611] = 8'b1101100;
DRAM[14612] = 8'b1101101;
DRAM[14613] = 8'b1101101;
DRAM[14614] = 8'b1101110;
DRAM[14615] = 8'b1101110;
DRAM[14616] = 8'b1110000;
DRAM[14617] = 8'b1110000;
DRAM[14618] = 8'b1110001;
DRAM[14619] = 8'b1110001;
DRAM[14620] = 8'b1110001;
DRAM[14621] = 8'b1110010;
DRAM[14622] = 8'b1110010;
DRAM[14623] = 8'b1110010;
DRAM[14624] = 8'b1110010;
DRAM[14625] = 8'b1110010;
DRAM[14626] = 8'b1110011;
DRAM[14627] = 8'b1110100;
DRAM[14628] = 8'b1110101;
DRAM[14629] = 8'b1110101;
DRAM[14630] = 8'b1110110;
DRAM[14631] = 8'b1110110;
DRAM[14632] = 8'b1101100;
DRAM[14633] = 8'b1110101;
DRAM[14634] = 8'b1110110;
DRAM[14635] = 8'b1111000;
DRAM[14636] = 8'b10000100;
DRAM[14637] = 8'b10000101;
DRAM[14638] = 8'b10000010;
DRAM[14639] = 8'b10000110;
DRAM[14640] = 8'b1111100;
DRAM[14641] = 8'b1111000;
DRAM[14642] = 8'b10001001;
DRAM[14643] = 8'b10110110;
DRAM[14644] = 8'b11100110;
DRAM[14645] = 8'b11111110;
DRAM[14646] = 8'b11111010;
DRAM[14647] = 8'b11110000;
DRAM[14648] = 8'b11111100;
DRAM[14649] = 8'b11111100;
DRAM[14650] = 8'b11111100;
DRAM[14651] = 8'b11111101;
DRAM[14652] = 8'b11111101;
DRAM[14653] = 8'b11111110;
DRAM[14654] = 8'b11111110;
DRAM[14655] = 8'b11111110;
DRAM[14656] = 8'b11111111;
DRAM[14657] = 8'b11111111;
DRAM[14658] = 8'b11111111;
DRAM[14659] = 8'b11111111;
DRAM[14660] = 8'b11111111;
DRAM[14661] = 8'b11111111;
DRAM[14662] = 8'b11111111;
DRAM[14663] = 8'b11111111;
DRAM[14664] = 8'b11111111;
DRAM[14665] = 8'b11111111;
DRAM[14666] = 8'b11111100;
DRAM[14667] = 8'b11111010;
DRAM[14668] = 8'b11111010;
DRAM[14669] = 8'b11111010;
DRAM[14670] = 8'b11111011;
DRAM[14671] = 8'b11111011;
DRAM[14672] = 8'b11110101;
DRAM[14673] = 8'b11111010;
DRAM[14674] = 8'b11111100;
DRAM[14675] = 8'b11111000;
DRAM[14676] = 8'b11110010;
DRAM[14677] = 8'b11101111;
DRAM[14678] = 8'b11110000;
DRAM[14679] = 8'b11110011;
DRAM[14680] = 8'b11101111;
DRAM[14681] = 8'b11110010;
DRAM[14682] = 8'b11110101;
DRAM[14683] = 8'b11110110;
DRAM[14684] = 8'b11111001;
DRAM[14685] = 8'b11111100;
DRAM[14686] = 8'b11111010;
DRAM[14687] = 8'b11110101;
DRAM[14688] = 8'b11110111;
DRAM[14689] = 8'b11111100;
DRAM[14690] = 8'b11111110;
DRAM[14691] = 8'b11111011;
DRAM[14692] = 8'b11111000;
DRAM[14693] = 8'b11111010;
DRAM[14694] = 8'b11111100;
DRAM[14695] = 8'b11111011;
DRAM[14696] = 8'b11110111;
DRAM[14697] = 8'b11111011;
DRAM[14698] = 8'b11111100;
DRAM[14699] = 8'b11111001;
DRAM[14700] = 8'b11110110;
DRAM[14701] = 8'b11110100;
DRAM[14702] = 8'b11110000;
DRAM[14703] = 8'b11101010;
DRAM[14704] = 8'b11101010;
DRAM[14705] = 8'b11110100;
DRAM[14706] = 8'b11111001;
DRAM[14707] = 8'b11110110;
DRAM[14708] = 8'b11110111;
DRAM[14709] = 8'b11111101;
DRAM[14710] = 8'b11111100;
DRAM[14711] = 8'b11110111;
DRAM[14712] = 8'b11110010;
DRAM[14713] = 8'b11110101;
DRAM[14714] = 8'b11110100;
DRAM[14715] = 8'b11110010;
DRAM[14716] = 8'b11110011;
DRAM[14717] = 8'b11110110;
DRAM[14718] = 8'b11110110;
DRAM[14719] = 8'b11110010;
DRAM[14720] = 8'b11110010;
DRAM[14721] = 8'b11110100;
DRAM[14722] = 8'b11110111;
DRAM[14723] = 8'b11111001;
DRAM[14724] = 8'b11111010;
DRAM[14725] = 8'b11111011;
DRAM[14726] = 8'b11111100;
DRAM[14727] = 8'b11111100;
DRAM[14728] = 8'b11110111;
DRAM[14729] = 8'b11111001;
DRAM[14730] = 8'b11111001;
DRAM[14731] = 8'b11110110;
DRAM[14732] = 8'b11110111;
DRAM[14733] = 8'b11111000;
DRAM[14734] = 8'b11110011;
DRAM[14735] = 8'b11101011;
DRAM[14736] = 8'b11110000;
DRAM[14737] = 8'b11101100;
DRAM[14738] = 8'b11110001;
DRAM[14739] = 8'b11110010;
DRAM[14740] = 8'b11101011;
DRAM[14741] = 8'b11101111;
DRAM[14742] = 8'b11110111;
DRAM[14743] = 8'b11110101;
DRAM[14744] = 8'b11111000;
DRAM[14745] = 8'b11101110;
DRAM[14746] = 8'b11101100;
DRAM[14747] = 8'b11110011;
DRAM[14748] = 8'b11110111;
DRAM[14749] = 8'b11110010;
DRAM[14750] = 8'b11110001;
DRAM[14751] = 8'b11110110;
DRAM[14752] = 8'b11110101;
DRAM[14753] = 8'b11110101;
DRAM[14754] = 8'b11110110;
DRAM[14755] = 8'b11111000;
DRAM[14756] = 8'b11111011;
DRAM[14757] = 8'b11111100;
DRAM[14758] = 8'b11111100;
DRAM[14759] = 8'b11111011;
DRAM[14760] = 8'b11111010;
DRAM[14761] = 8'b11111111;
DRAM[14762] = 8'b11111111;
DRAM[14763] = 8'b11111100;
DRAM[14764] = 8'b11111010;
DRAM[14765] = 8'b11111101;
DRAM[14766] = 8'b11111110;
DRAM[14767] = 8'b11111011;
DRAM[14768] = 8'b11110111;
DRAM[14769] = 8'b11111101;
DRAM[14770] = 8'b11111111;
DRAM[14771] = 8'b11111101;
DRAM[14772] = 8'b11111111;
DRAM[14773] = 8'b11111110;
DRAM[14774] = 8'b11101110;
DRAM[14775] = 8'b11011001;
DRAM[14776] = 8'b10110101;
DRAM[14777] = 8'b10110101;
DRAM[14778] = 8'b10110100;
DRAM[14779] = 8'b10110100;
DRAM[14780] = 8'b10111101;
DRAM[14781] = 8'b11010001;
DRAM[14782] = 8'b11101000;
DRAM[14783] = 8'b11110111;
DRAM[14784] = 8'b11111110;
DRAM[14785] = 8'b11110011;
DRAM[14786] = 8'b11111101;
DRAM[14787] = 8'b11111111;
DRAM[14788] = 8'b11111101;
DRAM[14789] = 8'b11111100;
DRAM[14790] = 8'b11111111;
DRAM[14791] = 8'b11111111;
DRAM[14792] = 8'b11111101;
DRAM[14793] = 8'b11111110;
DRAM[14794] = 8'b11111111;
DRAM[14795] = 8'b11111111;
DRAM[14796] = 8'b11111101;
DRAM[14797] = 8'b11111100;
DRAM[14798] = 8'b11111101;
DRAM[14799] = 8'b11111110;
DRAM[14800] = 8'b11111101;
DRAM[14801] = 8'b11111011;
DRAM[14802] = 8'b11111011;
DRAM[14803] = 8'b11111100;
DRAM[14804] = 8'b11111110;
DRAM[14805] = 8'b11111101;
DRAM[14806] = 8'b11111000;
DRAM[14807] = 8'b11110101;
DRAM[14808] = 8'b11101111;
DRAM[14809] = 8'b11001110;
DRAM[14810] = 8'b10100010;
DRAM[14811] = 8'b10000010;
DRAM[14812] = 8'b1110000;
DRAM[14813] = 8'b1100101;
DRAM[14814] = 8'b1011101;
DRAM[14815] = 8'b1011000;
DRAM[14816] = 8'b1100010;
DRAM[14817] = 8'b1100001;
DRAM[14818] = 8'b1011110;
DRAM[14819] = 8'b1011011;
DRAM[14820] = 8'b1011010;
DRAM[14821] = 8'b1011001;
DRAM[14822] = 8'b1011000;
DRAM[14823] = 8'b1010110;
DRAM[14824] = 8'b1010111;
DRAM[14825] = 8'b1011000;
DRAM[14826] = 8'b1011000;
DRAM[14827] = 8'b1011001;
DRAM[14828] = 8'b1011000;
DRAM[14829] = 8'b1010111;
DRAM[14830] = 8'b1010110;
DRAM[14831] = 8'b1010101;
DRAM[14832] = 8'b1010101;
DRAM[14833] = 8'b1010101;
DRAM[14834] = 8'b1010101;
DRAM[14835] = 8'b1010101;
DRAM[14836] = 8'b1010101;
DRAM[14837] = 8'b1010100;
DRAM[14838] = 8'b1010011;
DRAM[14839] = 8'b1010011;
DRAM[14840] = 8'b1010101;
DRAM[14841] = 8'b1010100;
DRAM[14842] = 8'b1010011;
DRAM[14843] = 8'b1010011;
DRAM[14844] = 8'b1010010;
DRAM[14845] = 8'b1010010;
DRAM[14846] = 8'b1010011;
DRAM[14847] = 8'b1010011;
DRAM[14848] = 8'b1100011;
DRAM[14849] = 8'b1100011;
DRAM[14850] = 8'b1100100;
DRAM[14851] = 8'b1100100;
DRAM[14852] = 8'b1100101;
DRAM[14853] = 8'b1100101;
DRAM[14854] = 8'b1100101;
DRAM[14855] = 8'b1100110;
DRAM[14856] = 8'b1100110;
DRAM[14857] = 8'b1100110;
DRAM[14858] = 8'b1100111;
DRAM[14859] = 8'b1101000;
DRAM[14860] = 8'b1101001;
DRAM[14861] = 8'b1101010;
DRAM[14862] = 8'b1101011;
DRAM[14863] = 8'b1101011;
DRAM[14864] = 8'b1101010;
DRAM[14865] = 8'b1101011;
DRAM[14866] = 8'b1101011;
DRAM[14867] = 8'b1101100;
DRAM[14868] = 8'b1101101;
DRAM[14869] = 8'b1101110;
DRAM[14870] = 8'b1101110;
DRAM[14871] = 8'b1101110;
DRAM[14872] = 8'b1110000;
DRAM[14873] = 8'b1110001;
DRAM[14874] = 8'b1110001;
DRAM[14875] = 8'b1110001;
DRAM[14876] = 8'b1110010;
DRAM[14877] = 8'b1110010;
DRAM[14878] = 8'b1110010;
DRAM[14879] = 8'b1110010;
DRAM[14880] = 8'b1110010;
DRAM[14881] = 8'b1110011;
DRAM[14882] = 8'b1110011;
DRAM[14883] = 8'b1110100;
DRAM[14884] = 8'b1110101;
DRAM[14885] = 8'b1110110;
DRAM[14886] = 8'b1110110;
DRAM[14887] = 8'b1110110;
DRAM[14888] = 8'b1111001;
DRAM[14889] = 8'b1111101;
DRAM[14890] = 8'b1111000;
DRAM[14891] = 8'b1111011;
DRAM[14892] = 8'b10000111;
DRAM[14893] = 8'b10001010;
DRAM[14894] = 8'b10001000;
DRAM[14895] = 8'b10001110;
DRAM[14896] = 8'b10011101;
DRAM[14897] = 8'b10100111;
DRAM[14898] = 8'b11000000;
DRAM[14899] = 8'b11100100;
DRAM[14900] = 8'b11111111;
DRAM[14901] = 8'b11111111;
DRAM[14902] = 8'b11111111;
DRAM[14903] = 8'b11111001;
DRAM[14904] = 8'b11111100;
DRAM[14905] = 8'b11111100;
DRAM[14906] = 8'b11111100;
DRAM[14907] = 8'b11111101;
DRAM[14908] = 8'b11111101;
DRAM[14909] = 8'b11111110;
DRAM[14910] = 8'b11111110;
DRAM[14911] = 8'b11111110;
DRAM[14912] = 8'b11111111;
DRAM[14913] = 8'b11111111;
DRAM[14914] = 8'b11111111;
DRAM[14915] = 8'b11111111;
DRAM[14916] = 8'b11111111;
DRAM[14917] = 8'b11111111;
DRAM[14918] = 8'b11111111;
DRAM[14919] = 8'b11111111;
DRAM[14920] = 8'b11111111;
DRAM[14921] = 8'b11111111;
DRAM[14922] = 8'b11111101;
DRAM[14923] = 8'b11111011;
DRAM[14924] = 8'b11111100;
DRAM[14925] = 8'b11111110;
DRAM[14926] = 8'b11111111;
DRAM[14927] = 8'b11111111;
DRAM[14928] = 8'b11111111;
DRAM[14929] = 8'b11111111;
DRAM[14930] = 8'b11110110;
DRAM[14931] = 8'b11100111;
DRAM[14932] = 8'b11011001;
DRAM[14933] = 8'b11010111;
DRAM[14934] = 8'b11100010;
DRAM[14935] = 8'b11101110;
DRAM[14936] = 8'b11101101;
DRAM[14937] = 8'b11110000;
DRAM[14938] = 8'b11110011;
DRAM[14939] = 8'b11110110;
DRAM[14940] = 8'b11111100;
DRAM[14941] = 8'b11111111;
DRAM[14942] = 8'b11111000;
DRAM[14943] = 8'b11101111;
DRAM[14944] = 8'b11110000;
DRAM[14945] = 8'b11110111;
DRAM[14946] = 8'b11111011;
DRAM[14947] = 8'b11111010;
DRAM[14948] = 8'b11111010;
DRAM[14949] = 8'b11111011;
DRAM[14950] = 8'b11111010;
DRAM[14951] = 8'b11110110;
DRAM[14952] = 8'b11111011;
DRAM[14953] = 8'b11111100;
DRAM[14954] = 8'b11111011;
DRAM[14955] = 8'b11111001;
DRAM[14956] = 8'b11111000;
DRAM[14957] = 8'b11110101;
DRAM[14958] = 8'b11101100;
DRAM[14959] = 8'b11100010;
DRAM[14960] = 8'b11100011;
DRAM[14961] = 8'b11101111;
DRAM[14962] = 8'b11110111;
DRAM[14963] = 8'b11110101;
DRAM[14964] = 8'b11110101;
DRAM[14965] = 8'b11111010;
DRAM[14966] = 8'b11111010;
DRAM[14967] = 8'b11110110;
DRAM[14968] = 8'b11110001;
DRAM[14969] = 8'b11110001;
DRAM[14970] = 8'b11101111;
DRAM[14971] = 8'b11101111;
DRAM[14972] = 8'b11110101;
DRAM[14973] = 8'b11111011;
DRAM[14974] = 8'b11111001;
DRAM[14975] = 8'b11110011;
DRAM[14976] = 8'b11101110;
DRAM[14977] = 8'b11110001;
DRAM[14978] = 8'b11110101;
DRAM[14979] = 8'b11111001;
DRAM[14980] = 8'b11111011;
DRAM[14981] = 8'b11111011;
DRAM[14982] = 8'b11111010;
DRAM[14983] = 8'b11111001;
DRAM[14984] = 8'b11110101;
DRAM[14985] = 8'b11110110;
DRAM[14986] = 8'b11110101;
DRAM[14987] = 8'b11110001;
DRAM[14988] = 8'b11110010;
DRAM[14989] = 8'b11110011;
DRAM[14990] = 8'b11110001;
DRAM[14991] = 8'b11101011;
DRAM[14992] = 8'b11110011;
DRAM[14993] = 8'b11101001;
DRAM[14994] = 8'b11101001;
DRAM[14995] = 8'b11101011;
DRAM[14996] = 8'b11101001;
DRAM[14997] = 8'b11110000;
DRAM[14998] = 8'b11110111;
DRAM[14999] = 8'b11110010;
DRAM[15000] = 8'b11110111;
DRAM[15001] = 8'b11101011;
DRAM[15002] = 8'b11100110;
DRAM[15003] = 8'b11101111;
DRAM[15004] = 8'b11110111;
DRAM[15005] = 8'b11110101;
DRAM[15006] = 8'b11110001;
DRAM[15007] = 8'b11110000;
DRAM[15008] = 8'b11101110;
DRAM[15009] = 8'b11110001;
DRAM[15010] = 8'b11110101;
DRAM[15011] = 8'b11111000;
DRAM[15012] = 8'b11111000;
DRAM[15013] = 8'b11111000;
DRAM[15014] = 8'b11111000;
DRAM[15015] = 8'b11111001;
DRAM[15016] = 8'b11111010;
DRAM[15017] = 8'b11111100;
DRAM[15018] = 8'b11111100;
DRAM[15019] = 8'b11111010;
DRAM[15020] = 8'b11111011;
DRAM[15021] = 8'b11111101;
DRAM[15022] = 8'b11111011;
DRAM[15023] = 8'b11110110;
DRAM[15024] = 8'b11101101;
DRAM[15025] = 8'b11110111;
DRAM[15026] = 8'b11111111;
DRAM[15027] = 8'b11111111;
DRAM[15028] = 8'b11110110;
DRAM[15029] = 8'b11011001;
DRAM[15030] = 8'b10101010;
DRAM[15031] = 8'b10000001;
DRAM[15032] = 8'b10101011;
DRAM[15033] = 8'b10100110;
DRAM[15034] = 8'b10100101;
DRAM[15035] = 8'b10101000;
DRAM[15036] = 8'b10101100;
DRAM[15037] = 8'b10111000;
DRAM[15038] = 8'b11010110;
DRAM[15039] = 8'b11110100;
DRAM[15040] = 8'b11111111;
DRAM[15041] = 8'b11111001;
DRAM[15042] = 8'b11111111;
DRAM[15043] = 8'b11111111;
DRAM[15044] = 8'b11111110;
DRAM[15045] = 8'b11111100;
DRAM[15046] = 8'b11111111;
DRAM[15047] = 8'b11111010;
DRAM[15048] = 8'b11111100;
DRAM[15049] = 8'b11111101;
DRAM[15050] = 8'b11111110;
DRAM[15051] = 8'b11111110;
DRAM[15052] = 8'b11111100;
DRAM[15053] = 8'b11111100;
DRAM[15054] = 8'b11111101;
DRAM[15055] = 8'b11111111;
DRAM[15056] = 8'b11111110;
DRAM[15057] = 8'b11111110;
DRAM[15058] = 8'b11111110;
DRAM[15059] = 8'b11111110;
DRAM[15060] = 8'b11111111;
DRAM[15061] = 8'b11111110;
DRAM[15062] = 8'b11111011;
DRAM[15063] = 8'b11111000;
DRAM[15064] = 8'b11111110;
DRAM[15065] = 8'b11110000;
DRAM[15066] = 8'b11001110;
DRAM[15067] = 8'b10011111;
DRAM[15068] = 8'b1111101;
DRAM[15069] = 8'b1101110;
DRAM[15070] = 8'b1100101;
DRAM[15071] = 8'b1011101;
DRAM[15072] = 8'b1011101;
DRAM[15073] = 8'b1011010;
DRAM[15074] = 8'b1011000;
DRAM[15075] = 8'b1011001;
DRAM[15076] = 8'b1011010;
DRAM[15077] = 8'b1011010;
DRAM[15078] = 8'b1011010;
DRAM[15079] = 8'b1011001;
DRAM[15080] = 8'b1011000;
DRAM[15081] = 8'b1011000;
DRAM[15082] = 8'b1011001;
DRAM[15083] = 8'b1011001;
DRAM[15084] = 8'b1011001;
DRAM[15085] = 8'b1011000;
DRAM[15086] = 8'b1010111;
DRAM[15087] = 8'b1010110;
DRAM[15088] = 8'b1010111;
DRAM[15089] = 8'b1010110;
DRAM[15090] = 8'b1010101;
DRAM[15091] = 8'b1010100;
DRAM[15092] = 8'b1010100;
DRAM[15093] = 8'b1010100;
DRAM[15094] = 8'b1010100;
DRAM[15095] = 8'b1010100;
DRAM[15096] = 8'b1010101;
DRAM[15097] = 8'b1010101;
DRAM[15098] = 8'b1010100;
DRAM[15099] = 8'b1010011;
DRAM[15100] = 8'b1010010;
DRAM[15101] = 8'b1010010;
DRAM[15102] = 8'b1010011;
DRAM[15103] = 8'b1010011;
DRAM[15104] = 8'b1100011;
DRAM[15105] = 8'b1100011;
DRAM[15106] = 8'b1100100;
DRAM[15107] = 8'b1100100;
DRAM[15108] = 8'b1100101;
DRAM[15109] = 8'b1100110;
DRAM[15110] = 8'b1100110;
DRAM[15111] = 8'b1100111;
DRAM[15112] = 8'b1100110;
DRAM[15113] = 8'b1100111;
DRAM[15114] = 8'b1100111;
DRAM[15115] = 8'b1101000;
DRAM[15116] = 8'b1101001;
DRAM[15117] = 8'b1101010;
DRAM[15118] = 8'b1101011;
DRAM[15119] = 8'b1101011;
DRAM[15120] = 8'b1101011;
DRAM[15121] = 8'b1101011;
DRAM[15122] = 8'b1101100;
DRAM[15123] = 8'b1101100;
DRAM[15124] = 8'b1101101;
DRAM[15125] = 8'b1101110;
DRAM[15126] = 8'b1101111;
DRAM[15127] = 8'b1101111;
DRAM[15128] = 8'b1110001;
DRAM[15129] = 8'b1110001;
DRAM[15130] = 8'b1110001;
DRAM[15131] = 8'b1110010;
DRAM[15132] = 8'b1110010;
DRAM[15133] = 8'b1110010;
DRAM[15134] = 8'b1110011;
DRAM[15135] = 8'b1110011;
DRAM[15136] = 8'b1110011;
DRAM[15137] = 8'b1110011;
DRAM[15138] = 8'b1110100;
DRAM[15139] = 8'b1110100;
DRAM[15140] = 8'b1110101;
DRAM[15141] = 8'b1110110;
DRAM[15142] = 8'b1110111;
DRAM[15143] = 8'b1110111;
DRAM[15144] = 8'b1111011;
DRAM[15145] = 8'b1111011;
DRAM[15146] = 8'b1110100;
DRAM[15147] = 8'b1110011;
DRAM[15148] = 8'b1111111;
DRAM[15149] = 8'b10000111;
DRAM[15150] = 8'b10010010;
DRAM[15151] = 8'b10100100;
DRAM[15152] = 8'b11001011;
DRAM[15153] = 8'b11011110;
DRAM[15154] = 8'b11110011;
DRAM[15155] = 8'b11111010;
DRAM[15156] = 8'b11110011;
DRAM[15157] = 8'b11101111;
DRAM[15158] = 8'b11111000;
DRAM[15159] = 8'b11111111;
DRAM[15160] = 8'b11111100;
DRAM[15161] = 8'b11111100;
DRAM[15162] = 8'b11111100;
DRAM[15163] = 8'b11111101;
DRAM[15164] = 8'b11111101;
DRAM[15165] = 8'b11111110;
DRAM[15166] = 8'b11111110;
DRAM[15167] = 8'b11111110;
DRAM[15168] = 8'b11111110;
DRAM[15169] = 8'b11111110;
DRAM[15170] = 8'b11111110;
DRAM[15171] = 8'b11111110;
DRAM[15172] = 8'b11111110;
DRAM[15173] = 8'b11111110;
DRAM[15174] = 8'b11111110;
DRAM[15175] = 8'b11111110;
DRAM[15176] = 8'b11111010;
DRAM[15177] = 8'b11111101;
DRAM[15178] = 8'b11111111;
DRAM[15179] = 8'b11111111;
DRAM[15180] = 8'b11111111;
DRAM[15181] = 8'b11111111;
DRAM[15182] = 8'b11111111;
DRAM[15183] = 8'b11111101;
DRAM[15184] = 8'b11101010;
DRAM[15185] = 8'b11100011;
DRAM[15186] = 8'b11011010;
DRAM[15187] = 8'b11010100;
DRAM[15188] = 8'b11010001;
DRAM[15189] = 8'b11010110;
DRAM[15190] = 8'b11100001;
DRAM[15191] = 8'b11101100;
DRAM[15192] = 8'b11101011;
DRAM[15193] = 8'b11110001;
DRAM[15194] = 8'b11110101;
DRAM[15195] = 8'b11110111;
DRAM[15196] = 8'b11111010;
DRAM[15197] = 8'b11111100;
DRAM[15198] = 8'b11111000;
DRAM[15199] = 8'b11110010;
DRAM[15200] = 8'b11101110;
DRAM[15201] = 8'b11110100;
DRAM[15202] = 8'b11110111;
DRAM[15203] = 8'b11110111;
DRAM[15204] = 8'b11111000;
DRAM[15205] = 8'b11111010;
DRAM[15206] = 8'b11111001;
DRAM[15207] = 8'b11110110;
DRAM[15208] = 8'b11111110;
DRAM[15209] = 8'b11111110;
DRAM[15210] = 8'b11111011;
DRAM[15211] = 8'b11111001;
DRAM[15212] = 8'b11111010;
DRAM[15213] = 8'b11110111;
DRAM[15214] = 8'b11101011;
DRAM[15215] = 8'b11011101;
DRAM[15216] = 8'b11100001;
DRAM[15217] = 8'b11101001;
DRAM[15218] = 8'b11101110;
DRAM[15219] = 8'b11101100;
DRAM[15220] = 8'b11101111;
DRAM[15221] = 8'b11110111;
DRAM[15222] = 8'b11111000;
DRAM[15223] = 8'b11110010;
DRAM[15224] = 8'b11101110;
DRAM[15225] = 8'b11110000;
DRAM[15226] = 8'b11101111;
DRAM[15227] = 8'b11101111;
DRAM[15228] = 8'b11110011;
DRAM[15229] = 8'b11111001;
DRAM[15230] = 8'b11111000;
DRAM[15231] = 8'b11110100;
DRAM[15232] = 8'b11101101;
DRAM[15233] = 8'b11110000;
DRAM[15234] = 8'b11110011;
DRAM[15235] = 8'b11111000;
DRAM[15236] = 8'b11111010;
DRAM[15237] = 8'b11111000;
DRAM[15238] = 8'b11110101;
DRAM[15239] = 8'b11110001;
DRAM[15240] = 8'b11110010;
DRAM[15241] = 8'b11110100;
DRAM[15242] = 8'b11110100;
DRAM[15243] = 8'b11110000;
DRAM[15244] = 8'b11101110;
DRAM[15245] = 8'b11101110;
DRAM[15246] = 8'b11101010;
DRAM[15247] = 8'b11100101;
DRAM[15248] = 8'b11110001;
DRAM[15249] = 8'b11101000;
DRAM[15250] = 8'b11101000;
DRAM[15251] = 8'b11101010;
DRAM[15252] = 8'b11101000;
DRAM[15253] = 8'b11101111;
DRAM[15254] = 8'b11110101;
DRAM[15255] = 8'b11110000;
DRAM[15256] = 8'b11110100;
DRAM[15257] = 8'b11101000;
DRAM[15258] = 8'b11100011;
DRAM[15259] = 8'b11101101;
DRAM[15260] = 8'b11111000;
DRAM[15261] = 8'b11111001;
DRAM[15262] = 8'b11110010;
DRAM[15263] = 8'b11101101;
DRAM[15264] = 8'b11101001;
DRAM[15265] = 8'b11101110;
DRAM[15266] = 8'b11110101;
DRAM[15267] = 8'b11111000;
DRAM[15268] = 8'b11110111;
DRAM[15269] = 8'b11110110;
DRAM[15270] = 8'b11110111;
DRAM[15271] = 8'b11111001;
DRAM[15272] = 8'b11111100;
DRAM[15273] = 8'b11111011;
DRAM[15274] = 8'b11111010;
DRAM[15275] = 8'b11111010;
DRAM[15276] = 8'b11111100;
DRAM[15277] = 8'b11111011;
DRAM[15278] = 8'b11110101;
DRAM[15279] = 8'b11110000;
DRAM[15280] = 8'b11110001;
DRAM[15281] = 8'b11110001;
DRAM[15282] = 8'b11101111;
DRAM[15283] = 8'b11110000;
DRAM[15284] = 8'b11111000;
DRAM[15285] = 8'b11111110;
DRAM[15286] = 8'b11111001;
DRAM[15287] = 8'b11101111;
DRAM[15288] = 8'b10111110;
DRAM[15289] = 8'b10101011;
DRAM[15290] = 8'b10011111;
DRAM[15291] = 8'b10100000;
DRAM[15292] = 8'b10011011;
DRAM[15293] = 8'b10011100;
DRAM[15294] = 8'b10110111;
DRAM[15295] = 8'b11011010;
DRAM[15296] = 8'b11111010;
DRAM[15297] = 8'b11111010;
DRAM[15298] = 8'b11111110;
DRAM[15299] = 8'b11111110;
DRAM[15300] = 8'b11111011;
DRAM[15301] = 8'b11111100;
DRAM[15302] = 8'b11111101;
DRAM[15303] = 8'b11111001;
DRAM[15304] = 8'b11111010;
DRAM[15305] = 8'b11111100;
DRAM[15306] = 8'b11111101;
DRAM[15307] = 8'b11111101;
DRAM[15308] = 8'b11111100;
DRAM[15309] = 8'b11111011;
DRAM[15310] = 8'b11111101;
DRAM[15311] = 8'b11111110;
DRAM[15312] = 8'b11111110;
DRAM[15313] = 8'b11111110;
DRAM[15314] = 8'b11111110;
DRAM[15315] = 8'b11111111;
DRAM[15316] = 8'b11111111;
DRAM[15317] = 8'b11111110;
DRAM[15318] = 8'b11111100;
DRAM[15319] = 8'b11111011;
DRAM[15320] = 8'b11111111;
DRAM[15321] = 8'b11111110;
DRAM[15322] = 8'b11101110;
DRAM[15323] = 8'b11001101;
DRAM[15324] = 8'b10101001;
DRAM[15325] = 8'b10001110;
DRAM[15326] = 8'b1111011;
DRAM[15327] = 8'b1101111;
DRAM[15328] = 8'b1100001;
DRAM[15329] = 8'b1011100;
DRAM[15330] = 8'b1011001;
DRAM[15331] = 8'b1011010;
DRAM[15332] = 8'b1011100;
DRAM[15333] = 8'b1011100;
DRAM[15334] = 8'b1011011;
DRAM[15335] = 8'b1011011;
DRAM[15336] = 8'b1011001;
DRAM[15337] = 8'b1011001;
DRAM[15338] = 8'b1011001;
DRAM[15339] = 8'b1011001;
DRAM[15340] = 8'b1011001;
DRAM[15341] = 8'b1011000;
DRAM[15342] = 8'b1011000;
DRAM[15343] = 8'b1010111;
DRAM[15344] = 8'b1011000;
DRAM[15345] = 8'b1010111;
DRAM[15346] = 8'b1010101;
DRAM[15347] = 8'b1010100;
DRAM[15348] = 8'b1010100;
DRAM[15349] = 8'b1010100;
DRAM[15350] = 8'b1010101;
DRAM[15351] = 8'b1010110;
DRAM[15352] = 8'b1010110;
DRAM[15353] = 8'b1010101;
DRAM[15354] = 8'b1010100;
DRAM[15355] = 8'b1010011;
DRAM[15356] = 8'b1010011;
DRAM[15357] = 8'b1010011;
DRAM[15358] = 8'b1010011;
DRAM[15359] = 8'b1010100;
DRAM[15360] = 8'b1100011;
DRAM[15361] = 8'b1100011;
DRAM[15362] = 8'b1100100;
DRAM[15363] = 8'b1100101;
DRAM[15364] = 8'b1100110;
DRAM[15365] = 8'b1100111;
DRAM[15366] = 8'b1100111;
DRAM[15367] = 8'b1101000;
DRAM[15368] = 8'b1100111;
DRAM[15369] = 8'b1101000;
DRAM[15370] = 8'b1101000;
DRAM[15371] = 8'b1101001;
DRAM[15372] = 8'b1101010;
DRAM[15373] = 8'b1101010;
DRAM[15374] = 8'b1101011;
DRAM[15375] = 8'b1101011;
DRAM[15376] = 8'b1101011;
DRAM[15377] = 8'b1101011;
DRAM[15378] = 8'b1101100;
DRAM[15379] = 8'b1101101;
DRAM[15380] = 8'b1101110;
DRAM[15381] = 8'b1101110;
DRAM[15382] = 8'b1101111;
DRAM[15383] = 8'b1101111;
DRAM[15384] = 8'b1110001;
DRAM[15385] = 8'b1110001;
DRAM[15386] = 8'b1110010;
DRAM[15387] = 8'b1110010;
DRAM[15388] = 8'b1110010;
DRAM[15389] = 8'b1110011;
DRAM[15390] = 8'b1110011;
DRAM[15391] = 8'b1110011;
DRAM[15392] = 8'b1110011;
DRAM[15393] = 8'b1110011;
DRAM[15394] = 8'b1110100;
DRAM[15395] = 8'b1110101;
DRAM[15396] = 8'b1110110;
DRAM[15397] = 8'b1110110;
DRAM[15398] = 8'b1110111;
DRAM[15399] = 8'b1110111;
DRAM[15400] = 8'b1110111;
DRAM[15401] = 8'b1111101;
DRAM[15402] = 8'b1111101;
DRAM[15403] = 8'b10000000;
DRAM[15404] = 8'b10001100;
DRAM[15405] = 8'b10011000;
DRAM[15406] = 8'b10110000;
DRAM[15407] = 8'b11001110;
DRAM[15408] = 8'b11011100;
DRAM[15409] = 8'b11101010;
DRAM[15410] = 8'b11111010;
DRAM[15411] = 8'b11111111;
DRAM[15412] = 8'b11111110;
DRAM[15413] = 8'b11111010;
DRAM[15414] = 8'b11111000;
DRAM[15415] = 8'b11111000;
DRAM[15416] = 8'b11111100;
DRAM[15417] = 8'b11111100;
DRAM[15418] = 8'b11111100;
DRAM[15419] = 8'b11111101;
DRAM[15420] = 8'b11111101;
DRAM[15421] = 8'b11111110;
DRAM[15422] = 8'b11111110;
DRAM[15423] = 8'b11111110;
DRAM[15424] = 8'b11111110;
DRAM[15425] = 8'b11111110;
DRAM[15426] = 8'b11111110;
DRAM[15427] = 8'b11111110;
DRAM[15428] = 8'b11111110;
DRAM[15429] = 8'b11111110;
DRAM[15430] = 8'b11111110;
DRAM[15431] = 8'b11111110;
DRAM[15432] = 8'b11111110;
DRAM[15433] = 8'b11111111;
DRAM[15434] = 8'b11111110;
DRAM[15435] = 8'b11111011;
DRAM[15436] = 8'b11111011;
DRAM[15437] = 8'b11111100;
DRAM[15438] = 8'b11110111;
DRAM[15439] = 8'b11101110;
DRAM[15440] = 8'b11011010;
DRAM[15441] = 8'b11010001;
DRAM[15442] = 8'b11001100;
DRAM[15443] = 8'b11010000;
DRAM[15444] = 8'b11010100;
DRAM[15445] = 8'b11010010;
DRAM[15446] = 8'b11001111;
DRAM[15447] = 8'b11001111;
DRAM[15448] = 8'b11101011;
DRAM[15449] = 8'b11110011;
DRAM[15450] = 8'b11111001;
DRAM[15451] = 8'b11110111;
DRAM[15452] = 8'b11110100;
DRAM[15453] = 8'b11110110;
DRAM[15454] = 8'b11111001;
DRAM[15455] = 8'b11111010;
DRAM[15456] = 8'b11110001;
DRAM[15457] = 8'b11110100;
DRAM[15458] = 8'b11110100;
DRAM[15459] = 8'b11110010;
DRAM[15460] = 8'b11110100;
DRAM[15461] = 8'b11111001;
DRAM[15462] = 8'b11111011;
DRAM[15463] = 8'b11111000;
DRAM[15464] = 8'b11111101;
DRAM[15465] = 8'b11111100;
DRAM[15466] = 8'b11111000;
DRAM[15467] = 8'b11110110;
DRAM[15468] = 8'b11111000;
DRAM[15469] = 8'b11110101;
DRAM[15470] = 8'b11101000;
DRAM[15471] = 8'b11011010;
DRAM[15472] = 8'b11100110;
DRAM[15473] = 8'b11101001;
DRAM[15474] = 8'b11100111;
DRAM[15475] = 8'b11100100;
DRAM[15476] = 8'b11101011;
DRAM[15477] = 8'b11110110;
DRAM[15478] = 8'b11111000;
DRAM[15479] = 8'b11110001;
DRAM[15480] = 8'b11101000;
DRAM[15481] = 8'b11101101;
DRAM[15482] = 8'b11101111;
DRAM[15483] = 8'b11101101;
DRAM[15484] = 8'b11101011;
DRAM[15485] = 8'b11101110;
DRAM[15486] = 8'b11110001;
DRAM[15487] = 8'b11110000;
DRAM[15488] = 8'b11101010;
DRAM[15489] = 8'b11101011;
DRAM[15490] = 8'b11101111;
DRAM[15491] = 8'b11110100;
DRAM[15492] = 8'b11110111;
DRAM[15493] = 8'b11110110;
DRAM[15494] = 8'b11110001;
DRAM[15495] = 8'b11101100;
DRAM[15496] = 8'b11101111;
DRAM[15497] = 8'b11110100;
DRAM[15498] = 8'b11110101;
DRAM[15499] = 8'b11110001;
DRAM[15500] = 8'b11101100;
DRAM[15501] = 8'b11101000;
DRAM[15502] = 8'b11100010;
DRAM[15503] = 8'b11011011;
DRAM[15504] = 8'b11101101;
DRAM[15505] = 8'b11100111;
DRAM[15506] = 8'b11101010;
DRAM[15507] = 8'b11101100;
DRAM[15508] = 8'b11101000;
DRAM[15509] = 8'b11101100;
DRAM[15510] = 8'b11110001;
DRAM[15511] = 8'b11101101;
DRAM[15512] = 8'b11110100;
DRAM[15513] = 8'b11101011;
DRAM[15514] = 8'b11100111;
DRAM[15515] = 8'b11101110;
DRAM[15516] = 8'b11110110;
DRAM[15517] = 8'b11110110;
DRAM[15518] = 8'b11101110;
DRAM[15519] = 8'b11100111;
DRAM[15520] = 8'b11100111;
DRAM[15521] = 8'b11101101;
DRAM[15522] = 8'b11110100;
DRAM[15523] = 8'b11110111;
DRAM[15524] = 8'b11110111;
DRAM[15525] = 8'b11110110;
DRAM[15526] = 8'b11111000;
DRAM[15527] = 8'b11111001;
DRAM[15528] = 8'b11111111;
DRAM[15529] = 8'b11111100;
DRAM[15530] = 8'b11111010;
DRAM[15531] = 8'b11111011;
DRAM[15532] = 8'b11111100;
DRAM[15533] = 8'b11111000;
DRAM[15534] = 8'b11110010;
DRAM[15535] = 8'b11101110;
DRAM[15536] = 8'b11101111;
DRAM[15537] = 8'b11110110;
DRAM[15538] = 8'b11111100;
DRAM[15539] = 8'b11111101;
DRAM[15540] = 8'b11111011;
DRAM[15541] = 8'b11110101;
DRAM[15542] = 8'b11101011;
DRAM[15543] = 8'b11100010;
DRAM[15544] = 8'b11001111;
DRAM[15545] = 8'b10101110;
DRAM[15546] = 8'b10010110;
DRAM[15547] = 8'b10010010;
DRAM[15548] = 8'b10001100;
DRAM[15549] = 8'b10000110;
DRAM[15550] = 8'b10011011;
DRAM[15551] = 8'b10111100;
DRAM[15552] = 8'b11101011;
DRAM[15553] = 8'b11110111;
DRAM[15554] = 8'b11111011;
DRAM[15555] = 8'b11111000;
DRAM[15556] = 8'b11111011;
DRAM[15557] = 8'b11111111;
DRAM[15558] = 8'b11111111;
DRAM[15559] = 8'b11111111;
DRAM[15560] = 8'b11111010;
DRAM[15561] = 8'b11111100;
DRAM[15562] = 8'b11111101;
DRAM[15563] = 8'b11111100;
DRAM[15564] = 8'b11111011;
DRAM[15565] = 8'b11111010;
DRAM[15566] = 8'b11111100;
DRAM[15567] = 8'b11111101;
DRAM[15568] = 8'b11111100;
DRAM[15569] = 8'b11111101;
DRAM[15570] = 8'b11111110;
DRAM[15571] = 8'b11111110;
DRAM[15572] = 8'b11111101;
DRAM[15573] = 8'b11111100;
DRAM[15574] = 8'b11111100;
DRAM[15575] = 8'b11111100;
DRAM[15576] = 8'b11111101;
DRAM[15577] = 8'b11111100;
DRAM[15578] = 8'b11111011;
DRAM[15579] = 8'b11110010;
DRAM[15580] = 8'b11010110;
DRAM[15581] = 8'b10101100;
DRAM[15582] = 8'b10000110;
DRAM[15583] = 8'b1110100;
DRAM[15584] = 8'b1110011;
DRAM[15585] = 8'b1101001;
DRAM[15586] = 8'b1100001;
DRAM[15587] = 8'b1100000;
DRAM[15588] = 8'b1100000;
DRAM[15589] = 8'b1011100;
DRAM[15590] = 8'b1011010;
DRAM[15591] = 8'b1011010;
DRAM[15592] = 8'b1011011;
DRAM[15593] = 8'b1011010;
DRAM[15594] = 8'b1011010;
DRAM[15595] = 8'b1011001;
DRAM[15596] = 8'b1011001;
DRAM[15597] = 8'b1011001;
DRAM[15598] = 8'b1011001;
DRAM[15599] = 8'b1011001;
DRAM[15600] = 8'b1011001;
DRAM[15601] = 8'b1011000;
DRAM[15602] = 8'b1010110;
DRAM[15603] = 8'b1010101;
DRAM[15604] = 8'b1010100;
DRAM[15605] = 8'b1010101;
DRAM[15606] = 8'b1010110;
DRAM[15607] = 8'b1010111;
DRAM[15608] = 8'b1010110;
DRAM[15609] = 8'b1010101;
DRAM[15610] = 8'b1010100;
DRAM[15611] = 8'b1010100;
DRAM[15612] = 8'b1010011;
DRAM[15613] = 8'b1010011;
DRAM[15614] = 8'b1010100;
DRAM[15615] = 8'b1010100;
DRAM[15616] = 8'b1100011;
DRAM[15617] = 8'b1100011;
DRAM[15618] = 8'b1100100;
DRAM[15619] = 8'b1100101;
DRAM[15620] = 8'b1100110;
DRAM[15621] = 8'b1100111;
DRAM[15622] = 8'b1101000;
DRAM[15623] = 8'b1101000;
DRAM[15624] = 8'b1101000;
DRAM[15625] = 8'b1101001;
DRAM[15626] = 8'b1101001;
DRAM[15627] = 8'b1101001;
DRAM[15628] = 8'b1101010;
DRAM[15629] = 8'b1101010;
DRAM[15630] = 8'b1101011;
DRAM[15631] = 8'b1101011;
DRAM[15632] = 8'b1101100;
DRAM[15633] = 8'b1101100;
DRAM[15634] = 8'b1101100;
DRAM[15635] = 8'b1101101;
DRAM[15636] = 8'b1101110;
DRAM[15637] = 8'b1101111;
DRAM[15638] = 8'b1101111;
DRAM[15639] = 8'b1110000;
DRAM[15640] = 8'b1110010;
DRAM[15641] = 8'b1110010;
DRAM[15642] = 8'b1110010;
DRAM[15643] = 8'b1110010;
DRAM[15644] = 8'b1110011;
DRAM[15645] = 8'b1110011;
DRAM[15646] = 8'b1110011;
DRAM[15647] = 8'b1110100;
DRAM[15648] = 8'b1110100;
DRAM[15649] = 8'b1110100;
DRAM[15650] = 8'b1110100;
DRAM[15651] = 8'b1110101;
DRAM[15652] = 8'b1110110;
DRAM[15653] = 8'b1110111;
DRAM[15654] = 8'b1110111;
DRAM[15655] = 8'b1111000;
DRAM[15656] = 8'b1110101;
DRAM[15657] = 8'b1111110;
DRAM[15658] = 8'b10000001;
DRAM[15659] = 8'b10000100;
DRAM[15660] = 8'b10001001;
DRAM[15661] = 8'b10001101;
DRAM[15662] = 8'b10100010;
DRAM[15663] = 8'b11000010;
DRAM[15664] = 8'b11100000;
DRAM[15665] = 8'b11101101;
DRAM[15666] = 8'b11111011;
DRAM[15667] = 8'b11111111;
DRAM[15668] = 8'b11111111;
DRAM[15669] = 8'b11111111;
DRAM[15670] = 8'b11111101;
DRAM[15671] = 8'b11111000;
DRAM[15672] = 8'b11111100;
DRAM[15673] = 8'b11111100;
DRAM[15674] = 8'b11111100;
DRAM[15675] = 8'b11111101;
DRAM[15676] = 8'b11111101;
DRAM[15677] = 8'b11111110;
DRAM[15678] = 8'b11111110;
DRAM[15679] = 8'b11111110;
DRAM[15680] = 8'b11111101;
DRAM[15681] = 8'b11111101;
DRAM[15682] = 8'b11111101;
DRAM[15683] = 8'b11111101;
DRAM[15684] = 8'b11111101;
DRAM[15685] = 8'b11111101;
DRAM[15686] = 8'b11111101;
DRAM[15687] = 8'b11111101;
DRAM[15688] = 8'b11111111;
DRAM[15689] = 8'b11111111;
DRAM[15690] = 8'b11111011;
DRAM[15691] = 8'b11110110;
DRAM[15692] = 8'b11111001;
DRAM[15693] = 8'b11111110;
DRAM[15694] = 8'b11110111;
DRAM[15695] = 8'b11101010;
DRAM[15696] = 8'b11011000;
DRAM[15697] = 8'b11001001;
DRAM[15698] = 8'b10111100;
DRAM[15699] = 8'b10111010;
DRAM[15700] = 8'b10111100;
DRAM[15701] = 8'b10111101;
DRAM[15702] = 8'b11000100;
DRAM[15703] = 8'b11001101;
DRAM[15704] = 8'b11101010;
DRAM[15705] = 8'b11110100;
DRAM[15706] = 8'b11111001;
DRAM[15707] = 8'b11110100;
DRAM[15708] = 8'b11101111;
DRAM[15709] = 8'b11110001;
DRAM[15710] = 8'b11111000;
DRAM[15711] = 8'b11111101;
DRAM[15712] = 8'b11110101;
DRAM[15713] = 8'b11110110;
DRAM[15714] = 8'b11110011;
DRAM[15715] = 8'b11101111;
DRAM[15716] = 8'b11110010;
DRAM[15717] = 8'b11111001;
DRAM[15718] = 8'b11111100;
DRAM[15719] = 8'b11111010;
DRAM[15720] = 8'b11111010;
DRAM[15721] = 8'b11111000;
DRAM[15722] = 8'b11110101;
DRAM[15723] = 8'b11110011;
DRAM[15724] = 8'b11110100;
DRAM[15725] = 8'b11110010;
DRAM[15726] = 8'b11100111;
DRAM[15727] = 8'b11011010;
DRAM[15728] = 8'b11101100;
DRAM[15729] = 8'b11101110;
DRAM[15730] = 8'b11101011;
DRAM[15731] = 8'b11100101;
DRAM[15732] = 8'b11101010;
DRAM[15733] = 8'b11110101;
DRAM[15734] = 8'b11111001;
DRAM[15735] = 8'b11110100;
DRAM[15736] = 8'b11100111;
DRAM[15737] = 8'b11101110;
DRAM[15738] = 8'b11110001;
DRAM[15739] = 8'b11101101;
DRAM[15740] = 8'b11101001;
DRAM[15741] = 8'b11101011;
DRAM[15742] = 8'b11101111;
DRAM[15743] = 8'b11110000;
DRAM[15744] = 8'b11100100;
DRAM[15745] = 8'b11100101;
DRAM[15746] = 8'b11101000;
DRAM[15747] = 8'b11101110;
DRAM[15748] = 8'b11110100;
DRAM[15749] = 8'b11110100;
DRAM[15750] = 8'b11110000;
DRAM[15751] = 8'b11101011;
DRAM[15752] = 8'b11101101;
DRAM[15753] = 8'b11110011;
DRAM[15754] = 8'b11110101;
DRAM[15755] = 8'b11110000;
DRAM[15756] = 8'b11101010;
DRAM[15757] = 8'b11100100;
DRAM[15758] = 8'b11011101;
DRAM[15759] = 8'b11010110;
DRAM[15760] = 8'b11101100;
DRAM[15761] = 8'b11100101;
DRAM[15762] = 8'b11101000;
DRAM[15763] = 8'b11101010;
DRAM[15764] = 8'b11100101;
DRAM[15765] = 8'b11101000;
DRAM[15766] = 8'b11101101;
DRAM[15767] = 8'b11100111;
DRAM[15768] = 8'b11110010;
DRAM[15769] = 8'b11101111;
DRAM[15770] = 8'b11101101;
DRAM[15771] = 8'b11101111;
DRAM[15772] = 8'b11110001;
DRAM[15773] = 8'b11101110;
DRAM[15774] = 8'b11100110;
DRAM[15775] = 8'b11100000;
DRAM[15776] = 8'b11101000;
DRAM[15777] = 8'b11101100;
DRAM[15778] = 8'b11110001;
DRAM[15779] = 8'b11110101;
DRAM[15780] = 8'b11110111;
DRAM[15781] = 8'b11111000;
DRAM[15782] = 8'b11111001;
DRAM[15783] = 8'b11111010;
DRAM[15784] = 8'b11111111;
DRAM[15785] = 8'b11111100;
DRAM[15786] = 8'b11111011;
DRAM[15787] = 8'b11111101;
DRAM[15788] = 8'b11111100;
DRAM[15789] = 8'b11110111;
DRAM[15790] = 8'b11110011;
DRAM[15791] = 8'b11110011;
DRAM[15792] = 8'b11111111;
DRAM[15793] = 8'b11111111;
DRAM[15794] = 8'b11111000;
DRAM[15795] = 8'b11101110;
DRAM[15796] = 8'b11101010;
DRAM[15797] = 8'b11101110;
DRAM[15798] = 8'b11111000;
DRAM[15799] = 8'b11111111;
DRAM[15800] = 8'b11001100;
DRAM[15801] = 8'b10100110;
DRAM[15802] = 8'b10001010;
DRAM[15803] = 8'b10001000;
DRAM[15804] = 8'b10001001;
DRAM[15805] = 8'b10001000;
DRAM[15806] = 8'b10011101;
DRAM[15807] = 8'b10111100;
DRAM[15808] = 8'b11100011;
DRAM[15809] = 8'b11111011;
DRAM[15810] = 8'b11111111;
DRAM[15811] = 8'b11111001;
DRAM[15812] = 8'b11111100;
DRAM[15813] = 8'b11111111;
DRAM[15814] = 8'b11111110;
DRAM[15815] = 8'b11111111;
DRAM[15816] = 8'b11111011;
DRAM[15817] = 8'b11111100;
DRAM[15818] = 8'b11111101;
DRAM[15819] = 8'b11111100;
DRAM[15820] = 8'b11111010;
DRAM[15821] = 8'b11111001;
DRAM[15822] = 8'b11111010;
DRAM[15823] = 8'b11111011;
DRAM[15824] = 8'b11111011;
DRAM[15825] = 8'b11111100;
DRAM[15826] = 8'b11111101;
DRAM[15827] = 8'b11111101;
DRAM[15828] = 8'b11111011;
DRAM[15829] = 8'b11111010;
DRAM[15830] = 8'b11111011;
DRAM[15831] = 8'b11111101;
DRAM[15832] = 8'b11111101;
DRAM[15833] = 8'b11111001;
DRAM[15834] = 8'b11111011;
DRAM[15835] = 8'b11111111;
DRAM[15836] = 8'b11101110;
DRAM[15837] = 8'b11000010;
DRAM[15838] = 8'b10010101;
DRAM[15839] = 8'b1111011;
DRAM[15840] = 8'b1110111;
DRAM[15841] = 8'b1101001;
DRAM[15842] = 8'b1011110;
DRAM[15843] = 8'b1011111;
DRAM[15844] = 8'b1100000;
DRAM[15845] = 8'b1011101;
DRAM[15846] = 8'b1011101;
DRAM[15847] = 8'b1100000;
DRAM[15848] = 8'b1011100;
DRAM[15849] = 8'b1011011;
DRAM[15850] = 8'b1011010;
DRAM[15851] = 8'b1011001;
DRAM[15852] = 8'b1011001;
DRAM[15853] = 8'b1011001;
DRAM[15854] = 8'b1011010;
DRAM[15855] = 8'b1011010;
DRAM[15856] = 8'b1011001;
DRAM[15857] = 8'b1011000;
DRAM[15858] = 8'b1010111;
DRAM[15859] = 8'b1010111;
DRAM[15860] = 8'b1010110;
DRAM[15861] = 8'b1010110;
DRAM[15862] = 8'b1010111;
DRAM[15863] = 8'b1010111;
DRAM[15864] = 8'b1010110;
DRAM[15865] = 8'b1010110;
DRAM[15866] = 8'b1010101;
DRAM[15867] = 8'b1010100;
DRAM[15868] = 8'b1010100;
DRAM[15869] = 8'b1010100;
DRAM[15870] = 8'b1010100;
DRAM[15871] = 8'b1010100;
DRAM[15872] = 8'b1100011;
DRAM[15873] = 8'b1100011;
DRAM[15874] = 8'b1100100;
DRAM[15875] = 8'b1100101;
DRAM[15876] = 8'b1100111;
DRAM[15877] = 8'b1101000;
DRAM[15878] = 8'b1101001;
DRAM[15879] = 8'b1101001;
DRAM[15880] = 8'b1101001;
DRAM[15881] = 8'b1101001;
DRAM[15882] = 8'b1101001;
DRAM[15883] = 8'b1101010;
DRAM[15884] = 8'b1101010;
DRAM[15885] = 8'b1101010;
DRAM[15886] = 8'b1101011;
DRAM[15887] = 8'b1101011;
DRAM[15888] = 8'b1101100;
DRAM[15889] = 8'b1101100;
DRAM[15890] = 8'b1101101;
DRAM[15891] = 8'b1101101;
DRAM[15892] = 8'b1101110;
DRAM[15893] = 8'b1101111;
DRAM[15894] = 8'b1110000;
DRAM[15895] = 8'b1110000;
DRAM[15896] = 8'b1110010;
DRAM[15897] = 8'b1110010;
DRAM[15898] = 8'b1110010;
DRAM[15899] = 8'b1110011;
DRAM[15900] = 8'b1110011;
DRAM[15901] = 8'b1110011;
DRAM[15902] = 8'b1110100;
DRAM[15903] = 8'b1110100;
DRAM[15904] = 8'b1110100;
DRAM[15905] = 8'b1110100;
DRAM[15906] = 8'b1110101;
DRAM[15907] = 8'b1110101;
DRAM[15908] = 8'b1110110;
DRAM[15909] = 8'b1110111;
DRAM[15910] = 8'b1111000;
DRAM[15911] = 8'b1111000;
DRAM[15912] = 8'b1110000;
DRAM[15913] = 8'b1110110;
DRAM[15914] = 8'b1110111;
DRAM[15915] = 8'b1111011;
DRAM[15916] = 8'b10000001;
DRAM[15917] = 8'b10000101;
DRAM[15918] = 8'b10011000;
DRAM[15919] = 8'b10111000;
DRAM[15920] = 8'b11101100;
DRAM[15921] = 8'b11111010;
DRAM[15922] = 8'b11111111;
DRAM[15923] = 8'b11111110;
DRAM[15924] = 8'b11110111;
DRAM[15925] = 8'b11111000;
DRAM[15926] = 8'b11111111;
DRAM[15927] = 8'b11111111;
DRAM[15928] = 8'b11111100;
DRAM[15929] = 8'b11111100;
DRAM[15930] = 8'b11111100;
DRAM[15931] = 8'b11111101;
DRAM[15932] = 8'b11111101;
DRAM[15933] = 8'b11111110;
DRAM[15934] = 8'b11111110;
DRAM[15935] = 8'b11111110;
DRAM[15936] = 8'b11111101;
DRAM[15937] = 8'b11111101;
DRAM[15938] = 8'b11111101;
DRAM[15939] = 8'b11111101;
DRAM[15940] = 8'b11111101;
DRAM[15941] = 8'b11111101;
DRAM[15942] = 8'b11111101;
DRAM[15943] = 8'b11111101;
DRAM[15944] = 8'b11111110;
DRAM[15945] = 8'b11111111;
DRAM[15946] = 8'b11111010;
DRAM[15947] = 8'b11110111;
DRAM[15948] = 8'b11111100;
DRAM[15949] = 8'b11111100;
DRAM[15950] = 8'b11101000;
DRAM[15951] = 8'b11010000;
DRAM[15952] = 8'b10101110;
DRAM[15953] = 8'b10100111;
DRAM[15954] = 8'b10100001;
DRAM[15955] = 8'b10011111;
DRAM[15956] = 8'b10011100;
DRAM[15957] = 8'b10100101;
DRAM[15958] = 8'b11000100;
DRAM[15959] = 8'b11100100;
DRAM[15960] = 8'b11101001;
DRAM[15961] = 8'b11110000;
DRAM[15962] = 8'b11110100;
DRAM[15963] = 8'b11110000;
DRAM[15964] = 8'b11101101;
DRAM[15965] = 8'b11110000;
DRAM[15966] = 8'b11110110;
DRAM[15967] = 8'b11111000;
DRAM[15968] = 8'b11111000;
DRAM[15969] = 8'b11110111;
DRAM[15970] = 8'b11110100;
DRAM[15971] = 8'b11110001;
DRAM[15972] = 8'b11110100;
DRAM[15973] = 8'b11111011;
DRAM[15974] = 8'b11111101;
DRAM[15975] = 8'b11111010;
DRAM[15976] = 8'b11111001;
DRAM[15977] = 8'b11111001;
DRAM[15978] = 8'b11110110;
DRAM[15979] = 8'b11110011;
DRAM[15980] = 8'b11110011;
DRAM[15981] = 8'b11110011;
DRAM[15982] = 8'b11101010;
DRAM[15983] = 8'b11100000;
DRAM[15984] = 8'b11101010;
DRAM[15985] = 8'b11110010;
DRAM[15986] = 8'b11110100;
DRAM[15987] = 8'b11101011;
DRAM[15988] = 8'b11101000;
DRAM[15989] = 8'b11101111;
DRAM[15990] = 8'b11110101;
DRAM[15991] = 8'b11110110;
DRAM[15992] = 8'b11101000;
DRAM[15993] = 8'b11101100;
DRAM[15994] = 8'b11101101;
DRAM[15995] = 8'b11101011;
DRAM[15996] = 8'b11101011;
DRAM[15997] = 8'b11101110;
DRAM[15998] = 8'b11101111;
DRAM[15999] = 8'b11101101;
DRAM[16000] = 8'b11100011;
DRAM[16001] = 8'b11100011;
DRAM[16002] = 8'b11100100;
DRAM[16003] = 8'b11101010;
DRAM[16004] = 8'b11101111;
DRAM[16005] = 8'b11110000;
DRAM[16006] = 8'b11101011;
DRAM[16007] = 8'b11100110;
DRAM[16008] = 8'b11101101;
DRAM[16009] = 8'b11110010;
DRAM[16010] = 8'b11110100;
DRAM[16011] = 8'b11101101;
DRAM[16012] = 8'b11100110;
DRAM[16013] = 8'b11100001;
DRAM[16014] = 8'b11011100;
DRAM[16015] = 8'b11010111;
DRAM[16016] = 8'b11110000;
DRAM[16017] = 8'b11100011;
DRAM[16018] = 8'b11100000;
DRAM[16019] = 8'b11100010;
DRAM[16020] = 8'b11100001;
DRAM[16021] = 8'b11100110;
DRAM[16022] = 8'b11101001;
DRAM[16023] = 8'b11100000;
DRAM[16024] = 8'b11100111;
DRAM[16025] = 8'b11101011;
DRAM[16026] = 8'b11101111;
DRAM[16027] = 8'b11101110;
DRAM[16028] = 8'b11101011;
DRAM[16029] = 8'b11100110;
DRAM[16030] = 8'b11100011;
DRAM[16031] = 8'b11100000;
DRAM[16032] = 8'b11101010;
DRAM[16033] = 8'b11101010;
DRAM[16034] = 8'b11101101;
DRAM[16035] = 8'b11110001;
DRAM[16036] = 8'b11110101;
DRAM[16037] = 8'b11111001;
DRAM[16038] = 8'b11111001;
DRAM[16039] = 8'b11111001;
DRAM[16040] = 8'b11111101;
DRAM[16041] = 8'b11111010;
DRAM[16042] = 8'b11111011;
DRAM[16043] = 8'b11111110;
DRAM[16044] = 8'b11111100;
DRAM[16045] = 8'b11110111;
DRAM[16046] = 8'b11111000;
DRAM[16047] = 8'b11111101;
DRAM[16048] = 8'b11110110;
DRAM[16049] = 8'b11111001;
DRAM[16050] = 8'b11111101;
DRAM[16051] = 8'b11111111;
DRAM[16052] = 8'b11111100;
DRAM[16053] = 8'b11110010;
DRAM[16054] = 8'b11101000;
DRAM[16055] = 8'b11100011;
DRAM[16056] = 8'b11010100;
DRAM[16057] = 8'b10110000;
DRAM[16058] = 8'b10010001;
DRAM[16059] = 8'b10001001;
DRAM[16060] = 8'b10000111;
DRAM[16061] = 8'b10001000;
DRAM[16062] = 8'b10011101;
DRAM[16063] = 8'b10111000;
DRAM[16064] = 8'b11001111;
DRAM[16065] = 8'b11110101;
DRAM[16066] = 8'b11111111;
DRAM[16067] = 8'b11111010;
DRAM[16068] = 8'b11111110;
DRAM[16069] = 8'b11111110;
DRAM[16070] = 8'b11111000;
DRAM[16071] = 8'b11111100;
DRAM[16072] = 8'b11111100;
DRAM[16073] = 8'b11111101;
DRAM[16074] = 8'b11111101;
DRAM[16075] = 8'b11111100;
DRAM[16076] = 8'b11111001;
DRAM[16077] = 8'b11110111;
DRAM[16078] = 8'b11111000;
DRAM[16079] = 8'b11111001;
DRAM[16080] = 8'b11111011;
DRAM[16081] = 8'b11111101;
DRAM[16082] = 8'b11111110;
DRAM[16083] = 8'b11111101;
DRAM[16084] = 8'b11111011;
DRAM[16085] = 8'b11111010;
DRAM[16086] = 8'b11111100;
DRAM[16087] = 8'b11111111;
DRAM[16088] = 8'b11111101;
DRAM[16089] = 8'b11111100;
DRAM[16090] = 8'b11111011;
DRAM[16091] = 8'b11111011;
DRAM[16092] = 8'b11111000;
DRAM[16093] = 8'b11100100;
DRAM[16094] = 8'b11000001;
DRAM[16095] = 8'b10100011;
DRAM[16096] = 8'b10000010;
DRAM[16097] = 8'b1101111;
DRAM[16098] = 8'b1100001;
DRAM[16099] = 8'b1100001;
DRAM[16100] = 8'b1100010;
DRAM[16101] = 8'b1011110;
DRAM[16102] = 8'b1011111;
DRAM[16103] = 8'b1100100;
DRAM[16104] = 8'b1011101;
DRAM[16105] = 8'b1011100;
DRAM[16106] = 8'b1011011;
DRAM[16107] = 8'b1011010;
DRAM[16108] = 8'b1011001;
DRAM[16109] = 8'b1011010;
DRAM[16110] = 8'b1011010;
DRAM[16111] = 8'b1011011;
DRAM[16112] = 8'b1011000;
DRAM[16113] = 8'b1011000;
DRAM[16114] = 8'b1011001;
DRAM[16115] = 8'b1011001;
DRAM[16116] = 8'b1011000;
DRAM[16117] = 8'b1010111;
DRAM[16118] = 8'b1010111;
DRAM[16119] = 8'b1010110;
DRAM[16120] = 8'b1010111;
DRAM[16121] = 8'b1010110;
DRAM[16122] = 8'b1010101;
DRAM[16123] = 8'b1010100;
DRAM[16124] = 8'b1010100;
DRAM[16125] = 8'b1010100;
DRAM[16126] = 8'b1010100;
DRAM[16127] = 8'b1010101;
DRAM[16128] = 8'b1100011;
DRAM[16129] = 8'b1100011;
DRAM[16130] = 8'b1100100;
DRAM[16131] = 8'b1100101;
DRAM[16132] = 8'b1100111;
DRAM[16133] = 8'b1101000;
DRAM[16134] = 8'b1101001;
DRAM[16135] = 8'b1101010;
DRAM[16136] = 8'b1101001;
DRAM[16137] = 8'b1101001;
DRAM[16138] = 8'b1101010;
DRAM[16139] = 8'b1101010;
DRAM[16140] = 8'b1101010;
DRAM[16141] = 8'b1101010;
DRAM[16142] = 8'b1101011;
DRAM[16143] = 8'b1101011;
DRAM[16144] = 8'b1101100;
DRAM[16145] = 8'b1101100;
DRAM[16146] = 8'b1101101;
DRAM[16147] = 8'b1101110;
DRAM[16148] = 8'b1101110;
DRAM[16149] = 8'b1101111;
DRAM[16150] = 8'b1110000;
DRAM[16151] = 8'b1110000;
DRAM[16152] = 8'b1110010;
DRAM[16153] = 8'b1110010;
DRAM[16154] = 8'b1110010;
DRAM[16155] = 8'b1110011;
DRAM[16156] = 8'b1110011;
DRAM[16157] = 8'b1110100;
DRAM[16158] = 8'b1110100;
DRAM[16159] = 8'b1110100;
DRAM[16160] = 8'b1110100;
DRAM[16161] = 8'b1110100;
DRAM[16162] = 8'b1110101;
DRAM[16163] = 8'b1110110;
DRAM[16164] = 8'b1110110;
DRAM[16165] = 8'b1110111;
DRAM[16166] = 8'b1111000;
DRAM[16167] = 8'b1111000;
DRAM[16168] = 8'b10000001;
DRAM[16169] = 8'b10000011;
DRAM[16170] = 8'b10000101;
DRAM[16171] = 8'b10010001;
DRAM[16172] = 8'b10100111;
DRAM[16173] = 8'b10111001;
DRAM[16174] = 8'b11011000;
DRAM[16175] = 8'b11111101;
DRAM[16176] = 8'b11110101;
DRAM[16177] = 8'b11111100;
DRAM[16178] = 8'b11111111;
DRAM[16179] = 8'b11111100;
DRAM[16180] = 8'b11111100;
DRAM[16181] = 8'b11111111;
DRAM[16182] = 8'b11111111;
DRAM[16183] = 8'b11111100;
DRAM[16184] = 8'b11111100;
DRAM[16185] = 8'b11111100;
DRAM[16186] = 8'b11111100;
DRAM[16187] = 8'b11111101;
DRAM[16188] = 8'b11111101;
DRAM[16189] = 8'b11111110;
DRAM[16190] = 8'b11111110;
DRAM[16191] = 8'b11111110;
DRAM[16192] = 8'b11111101;
DRAM[16193] = 8'b11111101;
DRAM[16194] = 8'b11111101;
DRAM[16195] = 8'b11111101;
DRAM[16196] = 8'b11111101;
DRAM[16197] = 8'b11111101;
DRAM[16198] = 8'b11111101;
DRAM[16199] = 8'b11111101;
DRAM[16200] = 8'b11111101;
DRAM[16201] = 8'b11111111;
DRAM[16202] = 8'b11111110;
DRAM[16203] = 8'b11111011;
DRAM[16204] = 8'b11111010;
DRAM[16205] = 8'b11101011;
DRAM[16206] = 8'b11000101;
DRAM[16207] = 8'b10011110;
DRAM[16208] = 8'b10010100;
DRAM[16209] = 8'b10011110;
DRAM[16210] = 8'b10101001;
DRAM[16211] = 8'b10100100;
DRAM[16212] = 8'b10001110;
DRAM[16213] = 8'b10000011;
DRAM[16214] = 8'b10011100;
DRAM[16215] = 8'b10111110;
DRAM[16216] = 8'b11101000;
DRAM[16217] = 8'b11101101;
DRAM[16218] = 8'b11101111;
DRAM[16219] = 8'b11101101;
DRAM[16220] = 8'b11101110;
DRAM[16221] = 8'b11110010;
DRAM[16222] = 8'b11110011;
DRAM[16223] = 8'b11110010;
DRAM[16224] = 8'b11111001;
DRAM[16225] = 8'b11111000;
DRAM[16226] = 8'b11110101;
DRAM[16227] = 8'b11110011;
DRAM[16228] = 8'b11110110;
DRAM[16229] = 8'b11111100;
DRAM[16230] = 8'b11111101;
DRAM[16231] = 8'b11111001;
DRAM[16232] = 8'b11111011;
DRAM[16233] = 8'b11111100;
DRAM[16234] = 8'b11111010;
DRAM[16235] = 8'b11110110;
DRAM[16236] = 8'b11110110;
DRAM[16237] = 8'b11110110;
DRAM[16238] = 8'b11110000;
DRAM[16239] = 8'b11101000;
DRAM[16240] = 8'b11100011;
DRAM[16241] = 8'b11110011;
DRAM[16242] = 8'b11111010;
DRAM[16243] = 8'b11101111;
DRAM[16244] = 8'b11100101;
DRAM[16245] = 8'b11100111;
DRAM[16246] = 8'b11110000;
DRAM[16247] = 8'b11110101;
DRAM[16248] = 8'b11100100;
DRAM[16249] = 8'b11100100;
DRAM[16250] = 8'b11100011;
DRAM[16251] = 8'b11100011;
DRAM[16252] = 8'b11100111;
DRAM[16253] = 8'b11101101;
DRAM[16254] = 8'b11101100;
DRAM[16255] = 8'b11100110;
DRAM[16256] = 8'b11100111;
DRAM[16257] = 8'b11100101;
DRAM[16258] = 8'b11100100;
DRAM[16259] = 8'b11101000;
DRAM[16260] = 8'b11101100;
DRAM[16261] = 8'b11101011;
DRAM[16262] = 8'b11100110;
DRAM[16263] = 8'b11100000;
DRAM[16264] = 8'b11101101;
DRAM[16265] = 8'b11110001;
DRAM[16266] = 8'b11110001;
DRAM[16267] = 8'b11101010;
DRAM[16268] = 8'b11100011;
DRAM[16269] = 8'b11100000;
DRAM[16270] = 8'b11011110;
DRAM[16271] = 8'b11011011;
DRAM[16272] = 8'b11110101;
DRAM[16273] = 8'b11100010;
DRAM[16274] = 8'b11011000;
DRAM[16275] = 8'b11011010;
DRAM[16276] = 8'b11011101;
DRAM[16277] = 8'b11100110;
DRAM[16278] = 8'b11100110;
DRAM[16279] = 8'b11011010;
DRAM[16280] = 8'b11011011;
DRAM[16281] = 8'b11100101;
DRAM[16282] = 8'b11101101;
DRAM[16283] = 8'b11101100;
DRAM[16284] = 8'b11100111;
DRAM[16285] = 8'b11100100;
DRAM[16286] = 8'b11100100;
DRAM[16287] = 8'b11100101;
DRAM[16288] = 8'b11101010;
DRAM[16289] = 8'b11101001;
DRAM[16290] = 8'b11101001;
DRAM[16291] = 8'b11101101;
DRAM[16292] = 8'b11110100;
DRAM[16293] = 8'b11111001;
DRAM[16294] = 8'b11111001;
DRAM[16295] = 8'b11111000;
DRAM[16296] = 8'b11111010;
DRAM[16297] = 8'b11111000;
DRAM[16298] = 8'b11111011;
DRAM[16299] = 8'b11111111;
DRAM[16300] = 8'b11111101;
DRAM[16301] = 8'b11111001;
DRAM[16302] = 8'b11111100;
DRAM[16303] = 8'b11111111;
DRAM[16304] = 8'b11111111;
DRAM[16305] = 8'b11111011;
DRAM[16306] = 8'b11111010;
DRAM[16307] = 8'b11111101;
DRAM[16308] = 8'b11111111;
DRAM[16309] = 8'b11111100;
DRAM[16310] = 8'b11110111;
DRAM[16311] = 8'b11110010;
DRAM[16312] = 8'b11101110;
DRAM[16313] = 8'b11001010;
DRAM[16314] = 8'b10100100;
DRAM[16315] = 8'b10001110;
DRAM[16316] = 8'b1111111;
DRAM[16317] = 8'b1110111;
DRAM[16318] = 8'b10000101;
DRAM[16319] = 8'b10011100;
DRAM[16320] = 8'b10101111;
DRAM[16321] = 8'b11100001;
DRAM[16322] = 8'b11111000;
DRAM[16323] = 8'b11110110;
DRAM[16324] = 8'b11111111;
DRAM[16325] = 8'b11111111;
DRAM[16326] = 8'b11111110;
DRAM[16327] = 8'b11111111;
DRAM[16328] = 8'b11111101;
DRAM[16329] = 8'b11111110;
DRAM[16330] = 8'b11111110;
DRAM[16331] = 8'b11111100;
DRAM[16332] = 8'b11111000;
DRAM[16333] = 8'b11110110;
DRAM[16334] = 8'b11110110;
DRAM[16335] = 8'b11110111;
DRAM[16336] = 8'b11111011;
DRAM[16337] = 8'b11111101;
DRAM[16338] = 8'b11111111;
DRAM[16339] = 8'b11111101;
DRAM[16340] = 8'b11111011;
DRAM[16341] = 8'b11111010;
DRAM[16342] = 8'b11111101;
DRAM[16343] = 8'b11111111;
DRAM[16344] = 8'b11111011;
DRAM[16345] = 8'b11111111;
DRAM[16346] = 8'b11111100;
DRAM[16347] = 8'b11110101;
DRAM[16348] = 8'b11111110;
DRAM[16349] = 8'b11111111;
DRAM[16350] = 8'b11110100;
DRAM[16351] = 8'b11010110;
DRAM[16352] = 8'b10100000;
DRAM[16353] = 8'b10001000;
DRAM[16354] = 8'b1110100;
DRAM[16355] = 8'b1101101;
DRAM[16356] = 8'b1101000;
DRAM[16357] = 8'b1011110;
DRAM[16358] = 8'b1011011;
DRAM[16359] = 8'b1011111;
DRAM[16360] = 8'b1011110;
DRAM[16361] = 8'b1011101;
DRAM[16362] = 8'b1011011;
DRAM[16363] = 8'b1011010;
DRAM[16364] = 8'b1011001;
DRAM[16365] = 8'b1011010;
DRAM[16366] = 8'b1011011;
DRAM[16367] = 8'b1011100;
DRAM[16368] = 8'b1010111;
DRAM[16369] = 8'b1011000;
DRAM[16370] = 8'b1011001;
DRAM[16371] = 8'b1011010;
DRAM[16372] = 8'b1011010;
DRAM[16373] = 8'b1011000;
DRAM[16374] = 8'b1010111;
DRAM[16375] = 8'b1010101;
DRAM[16376] = 8'b1010111;
DRAM[16377] = 8'b1010110;
DRAM[16378] = 8'b1010101;
DRAM[16379] = 8'b1010100;
DRAM[16380] = 8'b1010100;
DRAM[16381] = 8'b1010100;
DRAM[16382] = 8'b1010100;
DRAM[16383] = 8'b1010101;
DRAM[16384] = 8'b1100111;
DRAM[16385] = 8'b1100111;
DRAM[16386] = 8'b1100111;
DRAM[16387] = 8'b1101000;
DRAM[16388] = 8'b1101000;
DRAM[16389] = 8'b1101000;
DRAM[16390] = 8'b1101001;
DRAM[16391] = 8'b1101001;
DRAM[16392] = 8'b1101001;
DRAM[16393] = 8'b1101001;
DRAM[16394] = 8'b1101010;
DRAM[16395] = 8'b1101010;
DRAM[16396] = 8'b1101011;
DRAM[16397] = 8'b1101100;
DRAM[16398] = 8'b1101101;
DRAM[16399] = 8'b1101101;
DRAM[16400] = 8'b1101101;
DRAM[16401] = 8'b1101110;
DRAM[16402] = 8'b1101111;
DRAM[16403] = 8'b1110000;
DRAM[16404] = 8'b1110010;
DRAM[16405] = 8'b1110011;
DRAM[16406] = 8'b1110100;
DRAM[16407] = 8'b1110101;
DRAM[16408] = 8'b1110101;
DRAM[16409] = 8'b1110100;
DRAM[16410] = 8'b1110011;
DRAM[16411] = 8'b1110010;
DRAM[16412] = 8'b1110010;
DRAM[16413] = 8'b1110010;
DRAM[16414] = 8'b1110010;
DRAM[16415] = 8'b1110011;
DRAM[16416] = 8'b1110010;
DRAM[16417] = 8'b1110111;
DRAM[16418] = 8'b1110101;
DRAM[16419] = 8'b1110111;
DRAM[16420] = 8'b1111101;
DRAM[16421] = 8'b1110111;
DRAM[16422] = 8'b1110100;
DRAM[16423] = 8'b1111101;
DRAM[16424] = 8'b10010110;
DRAM[16425] = 8'b10010001;
DRAM[16426] = 8'b10100100;
DRAM[16427] = 8'b11001101;
DRAM[16428] = 8'b11101101;
DRAM[16429] = 8'b11110101;
DRAM[16430] = 8'b11111001;
DRAM[16431] = 8'b11111111;
DRAM[16432] = 8'b11111100;
DRAM[16433] = 8'b11111100;
DRAM[16434] = 8'b11111100;
DRAM[16435] = 8'b11111101;
DRAM[16436] = 8'b11111101;
DRAM[16437] = 8'b11111110;
DRAM[16438] = 8'b11111110;
DRAM[16439] = 8'b11111110;
DRAM[16440] = 8'b11111110;
DRAM[16441] = 8'b11111110;
DRAM[16442] = 8'b11111101;
DRAM[16443] = 8'b11111011;
DRAM[16444] = 8'b11111010;
DRAM[16445] = 8'b11111011;
DRAM[16446] = 8'b11111110;
DRAM[16447] = 8'b11111111;
DRAM[16448] = 8'b11111000;
DRAM[16449] = 8'b11111111;
DRAM[16450] = 8'b11111110;
DRAM[16451] = 8'b11111011;
DRAM[16452] = 8'b11111110;
DRAM[16453] = 8'b11111100;
DRAM[16454] = 8'b11111011;
DRAM[16455] = 8'b11111111;
DRAM[16456] = 8'b11111111;
DRAM[16457] = 8'b11110111;
DRAM[16458] = 8'b11101001;
DRAM[16459] = 8'b11111100;
DRAM[16460] = 8'b11111111;
DRAM[16461] = 8'b11010101;
DRAM[16462] = 8'b10011011;
DRAM[16463] = 8'b10011011;
DRAM[16464] = 8'b10100001;
DRAM[16465] = 8'b10101101;
DRAM[16466] = 8'b10010110;
DRAM[16467] = 8'b1111111;
DRAM[16468] = 8'b10010111;
DRAM[16469] = 8'b10111000;
DRAM[16470] = 8'b11000100;
DRAM[16471] = 8'b11001100;
DRAM[16472] = 8'b11010000;
DRAM[16473] = 8'b11011110;
DRAM[16474] = 8'b11101011;
DRAM[16475] = 8'b11101111;
DRAM[16476] = 8'b11110011;
DRAM[16477] = 8'b11110110;
DRAM[16478] = 8'b11101110;
DRAM[16479] = 8'b11100000;
DRAM[16480] = 8'b11110011;
DRAM[16481] = 8'b11110101;
DRAM[16482] = 8'b11110111;
DRAM[16483] = 8'b11111000;
DRAM[16484] = 8'b11110110;
DRAM[16485] = 8'b11110100;
DRAM[16486] = 8'b11110100;
DRAM[16487] = 8'b11110011;
DRAM[16488] = 8'b11111111;
DRAM[16489] = 8'b11111011;
DRAM[16490] = 8'b11110101;
DRAM[16491] = 8'b11110101;
DRAM[16492] = 8'b11111001;
DRAM[16493] = 8'b11111100;
DRAM[16494] = 8'b11111010;
DRAM[16495] = 8'b11110110;
DRAM[16496] = 8'b11011011;
DRAM[16497] = 8'b11100110;
DRAM[16498] = 8'b11101011;
DRAM[16499] = 8'b11100110;
DRAM[16500] = 8'b11110110;
DRAM[16501] = 8'b11110001;
DRAM[16502] = 8'b11011100;
DRAM[16503] = 8'b11110010;
DRAM[16504] = 8'b11101110;
DRAM[16505] = 8'b11011010;
DRAM[16506] = 8'b11011101;
DRAM[16507] = 8'b11100111;
DRAM[16508] = 8'b11100100;
DRAM[16509] = 8'b11101011;
DRAM[16510] = 8'b11101101;
DRAM[16511] = 8'b11011011;
DRAM[16512] = 8'b11101000;
DRAM[16513] = 8'b11011110;
DRAM[16514] = 8'b11011011;
DRAM[16515] = 8'b11011101;
DRAM[16516] = 8'b11011110;
DRAM[16517] = 8'b11101001;
DRAM[16518] = 8'b11110000;
DRAM[16519] = 8'b11101001;
DRAM[16520] = 8'b11101000;
DRAM[16521] = 8'b11110000;
DRAM[16522] = 8'b11110101;
DRAM[16523] = 8'b11011100;
DRAM[16524] = 8'b11110001;
DRAM[16525] = 8'b11100000;
DRAM[16526] = 8'b11010001;
DRAM[16527] = 8'b11100111;
DRAM[16528] = 8'b11110010;
DRAM[16529] = 8'b11100110;
DRAM[16530] = 8'b11100001;
DRAM[16531] = 8'b11100000;
DRAM[16532] = 8'b11011101;
DRAM[16533] = 8'b11011111;
DRAM[16534] = 8'b11011111;
DRAM[16535] = 8'b11010110;
DRAM[16536] = 8'b11100100;
DRAM[16537] = 8'b11101001;
DRAM[16538] = 8'b11011000;
DRAM[16539] = 8'b11100011;
DRAM[16540] = 8'b11100011;
DRAM[16541] = 8'b11011011;
DRAM[16542] = 8'b11101111;
DRAM[16543] = 8'b11101101;
DRAM[16544] = 8'b11100111;
DRAM[16545] = 8'b11100001;
DRAM[16546] = 8'b11101011;
DRAM[16547] = 8'b11101110;
DRAM[16548] = 8'b11100101;
DRAM[16549] = 8'b11101110;
DRAM[16550] = 8'b11111000;
DRAM[16551] = 8'b11101101;
DRAM[16552] = 8'b11110010;
DRAM[16553] = 8'b11110100;
DRAM[16554] = 8'b11110111;
DRAM[16555] = 8'b11111001;
DRAM[16556] = 8'b11111011;
DRAM[16557] = 8'b11111011;
DRAM[16558] = 8'b11111010;
DRAM[16559] = 8'b11111001;
DRAM[16560] = 8'b11110101;
DRAM[16561] = 8'b11110000;
DRAM[16562] = 8'b11101100;
DRAM[16563] = 8'b11101110;
DRAM[16564] = 8'b11110011;
DRAM[16565] = 8'b11110101;
DRAM[16566] = 8'b11110001;
DRAM[16567] = 8'b11101100;
DRAM[16568] = 8'b11010101;
DRAM[16569] = 8'b11001110;
DRAM[16570] = 8'b11011101;
DRAM[16571] = 8'b11001000;
DRAM[16572] = 8'b10101001;
DRAM[16573] = 8'b10101101;
DRAM[16574] = 8'b10101011;
DRAM[16575] = 8'b10100011;
DRAM[16576] = 8'b10100100;
DRAM[16577] = 8'b11010100;
DRAM[16578] = 8'b11111010;
DRAM[16579] = 8'b11110001;
DRAM[16580] = 8'b11111111;
DRAM[16581] = 8'b11111010;
DRAM[16582] = 8'b11111110;
DRAM[16583] = 8'b11111111;
DRAM[16584] = 8'b11111110;
DRAM[16585] = 8'b11111110;
DRAM[16586] = 8'b11111100;
DRAM[16587] = 8'b11111011;
DRAM[16588] = 8'b11111101;
DRAM[16589] = 8'b11111010;
DRAM[16590] = 8'b11101110;
DRAM[16591] = 8'b11100000;
DRAM[16592] = 8'b11100111;
DRAM[16593] = 8'b11110000;
DRAM[16594] = 8'b11111100;
DRAM[16595] = 8'b11111111;
DRAM[16596] = 8'b11111111;
DRAM[16597] = 8'b11111100;
DRAM[16598] = 8'b11111011;
DRAM[16599] = 8'b11111100;
DRAM[16600] = 8'b11111100;
DRAM[16601] = 8'b11111100;
DRAM[16602] = 8'b11111101;
DRAM[16603] = 8'b11111100;
DRAM[16604] = 8'b11111011;
DRAM[16605] = 8'b11111000;
DRAM[16606] = 8'b11110110;
DRAM[16607] = 8'b11110100;
DRAM[16608] = 8'b11000100;
DRAM[16609] = 8'b10011110;
DRAM[16610] = 8'b10001010;
DRAM[16611] = 8'b10000011;
DRAM[16612] = 8'b1110010;
DRAM[16613] = 8'b1101011;
DRAM[16614] = 8'b1100110;
DRAM[16615] = 8'b1010110;
DRAM[16616] = 8'b1011010;
DRAM[16617] = 8'b1011111;
DRAM[16618] = 8'b1100000;
DRAM[16619] = 8'b1011010;
DRAM[16620] = 8'b1011001;
DRAM[16621] = 8'b1011101;
DRAM[16622] = 8'b1011101;
DRAM[16623] = 8'b1011010;
DRAM[16624] = 8'b1011001;
DRAM[16625] = 8'b1011001;
DRAM[16626] = 8'b1011000;
DRAM[16627] = 8'b1011000;
DRAM[16628] = 8'b1011000;
DRAM[16629] = 8'b1010111;
DRAM[16630] = 8'b1010111;
DRAM[16631] = 8'b1010111;
DRAM[16632] = 8'b1011000;
DRAM[16633] = 8'b1010111;
DRAM[16634] = 8'b1010110;
DRAM[16635] = 8'b1010101;
DRAM[16636] = 8'b1010101;
DRAM[16637] = 8'b1010101;
DRAM[16638] = 8'b1010101;
DRAM[16639] = 8'b1010110;
DRAM[16640] = 8'b1100111;
DRAM[16641] = 8'b1100111;
DRAM[16642] = 8'b1101000;
DRAM[16643] = 8'b1101000;
DRAM[16644] = 8'b1101000;
DRAM[16645] = 8'b1101001;
DRAM[16646] = 8'b1101001;
DRAM[16647] = 8'b1101001;
DRAM[16648] = 8'b1101001;
DRAM[16649] = 8'b1101001;
DRAM[16650] = 8'b1101010;
DRAM[16651] = 8'b1101011;
DRAM[16652] = 8'b1101100;
DRAM[16653] = 8'b1101100;
DRAM[16654] = 8'b1101101;
DRAM[16655] = 8'b1101101;
DRAM[16656] = 8'b1101110;
DRAM[16657] = 8'b1101110;
DRAM[16658] = 8'b1101111;
DRAM[16659] = 8'b1110000;
DRAM[16660] = 8'b1110001;
DRAM[16661] = 8'b1110010;
DRAM[16662] = 8'b1110011;
DRAM[16663] = 8'b1110011;
DRAM[16664] = 8'b1110011;
DRAM[16665] = 8'b1110010;
DRAM[16666] = 8'b1110010;
DRAM[16667] = 8'b1110010;
DRAM[16668] = 8'b1110011;
DRAM[16669] = 8'b1110100;
DRAM[16670] = 8'b1110101;
DRAM[16671] = 8'b1110101;
DRAM[16672] = 8'b1110101;
DRAM[16673] = 8'b1110110;
DRAM[16674] = 8'b1110001;
DRAM[16675] = 8'b1110010;
DRAM[16676] = 8'b1111010;
DRAM[16677] = 8'b1111000;
DRAM[16678] = 8'b1110111;
DRAM[16679] = 8'b10000001;
DRAM[16680] = 8'b1111110;
DRAM[16681] = 8'b10001110;
DRAM[16682] = 8'b10110011;
DRAM[16683] = 8'b11011111;
DRAM[16684] = 8'b11111001;
DRAM[16685] = 8'b11111100;
DRAM[16686] = 8'b11111011;
DRAM[16687] = 8'b11111101;
DRAM[16688] = 8'b11111011;
DRAM[16689] = 8'b11111100;
DRAM[16690] = 8'b11111101;
DRAM[16691] = 8'b11111110;
DRAM[16692] = 8'b11111110;
DRAM[16693] = 8'b11111110;
DRAM[16694] = 8'b11111110;
DRAM[16695] = 8'b11111110;
DRAM[16696] = 8'b11111101;
DRAM[16697] = 8'b11111100;
DRAM[16698] = 8'b11111011;
DRAM[16699] = 8'b11111010;
DRAM[16700] = 8'b11111010;
DRAM[16701] = 8'b11111011;
DRAM[16702] = 8'b11111110;
DRAM[16703] = 8'b11111111;
DRAM[16704] = 8'b11111011;
DRAM[16705] = 8'b11111111;
DRAM[16706] = 8'b11111011;
DRAM[16707] = 8'b11111010;
DRAM[16708] = 8'b11111111;
DRAM[16709] = 8'b11111110;
DRAM[16710] = 8'b11111010;
DRAM[16711] = 8'b11111101;
DRAM[16712] = 8'b11101111;
DRAM[16713] = 8'b11110111;
DRAM[16714] = 8'b11110000;
DRAM[16715] = 8'b11101011;
DRAM[16716] = 8'b11101111;
DRAM[16717] = 8'b11011100;
DRAM[16718] = 8'b10111111;
DRAM[16719] = 8'b10111001;
DRAM[16720] = 8'b10010000;
DRAM[16721] = 8'b10010111;
DRAM[16722] = 8'b1111101;
DRAM[16723] = 8'b1100010;
DRAM[16724] = 8'b1110110;
DRAM[16725] = 8'b10011110;
DRAM[16726] = 8'b10111110;
DRAM[16727] = 8'b11010111;
DRAM[16728] = 8'b11011111;
DRAM[16729] = 8'b11011001;
DRAM[16730] = 8'b11010110;
DRAM[16731] = 8'b11011101;
DRAM[16732] = 8'b11101110;
DRAM[16733] = 8'b11111000;
DRAM[16734] = 8'b11110000;
DRAM[16735] = 8'b11100011;
DRAM[16736] = 8'b11101110;
DRAM[16737] = 8'b11110001;
DRAM[16738] = 8'b11110011;
DRAM[16739] = 8'b11110001;
DRAM[16740] = 8'b11101111;
DRAM[16741] = 8'b11110000;
DRAM[16742] = 8'b11110110;
DRAM[16743] = 8'b11111011;
DRAM[16744] = 8'b11110011;
DRAM[16745] = 8'b11110100;
DRAM[16746] = 8'b11110111;
DRAM[16747] = 8'b11111001;
DRAM[16748] = 8'b11111010;
DRAM[16749] = 8'b11111000;
DRAM[16750] = 8'b11110100;
DRAM[16751] = 8'b11110001;
DRAM[16752] = 8'b11101100;
DRAM[16753] = 8'b11100010;
DRAM[16754] = 8'b11110000;
DRAM[16755] = 8'b11101110;
DRAM[16756] = 8'b11100111;
DRAM[16757] = 8'b11101000;
DRAM[16758] = 8'b11100000;
DRAM[16759] = 8'b11100101;
DRAM[16760] = 8'b11101010;
DRAM[16761] = 8'b11011000;
DRAM[16762] = 8'b11011001;
DRAM[16763] = 8'b11100001;
DRAM[16764] = 8'b11011111;
DRAM[16765] = 8'b11100111;
DRAM[16766] = 8'b11101111;
DRAM[16767] = 8'b11100101;
DRAM[16768] = 8'b11101011;
DRAM[16769] = 8'b11100101;
DRAM[16770] = 8'b11100110;
DRAM[16771] = 8'b11100101;
DRAM[16772] = 8'b11100000;
DRAM[16773] = 8'b11100101;
DRAM[16774] = 8'b11101101;
DRAM[16775] = 8'b11101010;
DRAM[16776] = 8'b11100010;
DRAM[16777] = 8'b11101001;
DRAM[16778] = 8'b11110001;
DRAM[16779] = 8'b11011011;
DRAM[16780] = 8'b11110000;
DRAM[16781] = 8'b11100000;
DRAM[16782] = 8'b11010110;
DRAM[16783] = 8'b11101100;
DRAM[16784] = 8'b11100111;
DRAM[16785] = 8'b11100000;
DRAM[16786] = 8'b11011100;
DRAM[16787] = 8'b11100000;
DRAM[16788] = 8'b11100110;
DRAM[16789] = 8'b11100101;
DRAM[16790] = 8'b11011010;
DRAM[16791] = 8'b11001111;
DRAM[16792] = 8'b11100000;
DRAM[16793] = 8'b11100110;
DRAM[16794] = 8'b11011000;
DRAM[16795] = 8'b11011111;
DRAM[16796] = 8'b11100000;
DRAM[16797] = 8'b11011100;
DRAM[16798] = 8'b11101110;
DRAM[16799] = 8'b11101010;
DRAM[16800] = 8'b11100011;
DRAM[16801] = 8'b11100101;
DRAM[16802] = 8'b11101100;
DRAM[16803] = 8'b11101011;
DRAM[16804] = 8'b11100110;
DRAM[16805] = 8'b11101100;
DRAM[16806] = 8'b11110011;
DRAM[16807] = 8'b11110000;
DRAM[16808] = 8'b11110110;
DRAM[16809] = 8'b11110111;
DRAM[16810] = 8'b11111010;
DRAM[16811] = 8'b11111101;
DRAM[16812] = 8'b11111110;
DRAM[16813] = 8'b11111110;
DRAM[16814] = 8'b11111101;
DRAM[16815] = 8'b11111100;
DRAM[16816] = 8'b11111011;
DRAM[16817] = 8'b11111010;
DRAM[16818] = 8'b11111001;
DRAM[16819] = 8'b11111000;
DRAM[16820] = 8'b11111001;
DRAM[16821] = 8'b11111000;
DRAM[16822] = 8'b11110111;
DRAM[16823] = 8'b11110111;
DRAM[16824] = 8'b11111000;
DRAM[16825] = 8'b11101110;
DRAM[16826] = 8'b11110011;
DRAM[16827] = 8'b11001110;
DRAM[16828] = 8'b10011010;
DRAM[16829] = 8'b10001000;
DRAM[16830] = 8'b1111111;
DRAM[16831] = 8'b1111100;
DRAM[16832] = 8'b10011010;
DRAM[16833] = 8'b11000010;
DRAM[16834] = 8'b11101001;
DRAM[16835] = 8'b11110001;
DRAM[16836] = 8'b11111101;
DRAM[16837] = 8'b11111001;
DRAM[16838] = 8'b11111010;
DRAM[16839] = 8'b11111010;
DRAM[16840] = 8'b11111011;
DRAM[16841] = 8'b11111011;
DRAM[16842] = 8'b11111010;
DRAM[16843] = 8'b11111010;
DRAM[16844] = 8'b11111101;
DRAM[16845] = 8'b11111100;
DRAM[16846] = 8'b11110001;
DRAM[16847] = 8'b11100101;
DRAM[16848] = 8'b11011100;
DRAM[16849] = 8'b11100001;
DRAM[16850] = 8'b11101011;
DRAM[16851] = 8'b11110100;
DRAM[16852] = 8'b11111100;
DRAM[16853] = 8'b11111111;
DRAM[16854] = 8'b11111111;
DRAM[16855] = 8'b11111111;
DRAM[16856] = 8'b11111010;
DRAM[16857] = 8'b11111011;
DRAM[16858] = 8'b11111101;
DRAM[16859] = 8'b11111110;
DRAM[16860] = 8'b11111110;
DRAM[16861] = 8'b11111101;
DRAM[16862] = 8'b11111100;
DRAM[16863] = 8'b11111011;
DRAM[16864] = 8'b11110110;
DRAM[16865] = 8'b11011101;
DRAM[16866] = 8'b10111011;
DRAM[16867] = 8'b10010101;
DRAM[16868] = 8'b1110010;
DRAM[16869] = 8'b1100110;
DRAM[16870] = 8'b1101000;
DRAM[16871] = 8'b1100110;
DRAM[16872] = 8'b1011011;
DRAM[16873] = 8'b1011111;
DRAM[16874] = 8'b1011111;
DRAM[16875] = 8'b1011010;
DRAM[16876] = 8'b1011000;
DRAM[16877] = 8'b1011100;
DRAM[16878] = 8'b1011100;
DRAM[16879] = 8'b1011001;
DRAM[16880] = 8'b1011001;
DRAM[16881] = 8'b1011001;
DRAM[16882] = 8'b1011001;
DRAM[16883] = 8'b1011001;
DRAM[16884] = 8'b1011000;
DRAM[16885] = 8'b1011000;
DRAM[16886] = 8'b1010111;
DRAM[16887] = 8'b1010111;
DRAM[16888] = 8'b1011000;
DRAM[16889] = 8'b1010111;
DRAM[16890] = 8'b1010111;
DRAM[16891] = 8'b1010110;
DRAM[16892] = 8'b1010101;
DRAM[16893] = 8'b1010101;
DRAM[16894] = 8'b1010110;
DRAM[16895] = 8'b1010110;
DRAM[16896] = 8'b1101000;
DRAM[16897] = 8'b1101000;
DRAM[16898] = 8'b1101000;
DRAM[16899] = 8'b1101001;
DRAM[16900] = 8'b1101001;
DRAM[16901] = 8'b1101001;
DRAM[16902] = 8'b1101010;
DRAM[16903] = 8'b1101010;
DRAM[16904] = 8'b1101010;
DRAM[16905] = 8'b1101010;
DRAM[16906] = 8'b1101011;
DRAM[16907] = 8'b1101011;
DRAM[16908] = 8'b1101100;
DRAM[16909] = 8'b1101101;
DRAM[16910] = 8'b1101110;
DRAM[16911] = 8'b1101110;
DRAM[16912] = 8'b1101111;
DRAM[16913] = 8'b1101111;
DRAM[16914] = 8'b1110000;
DRAM[16915] = 8'b1110000;
DRAM[16916] = 8'b1110001;
DRAM[16917] = 8'b1110001;
DRAM[16918] = 8'b1110010;
DRAM[16919] = 8'b1110010;
DRAM[16920] = 8'b1110001;
DRAM[16921] = 8'b1110001;
DRAM[16922] = 8'b1110010;
DRAM[16923] = 8'b1110010;
DRAM[16924] = 8'b1110100;
DRAM[16925] = 8'b1110101;
DRAM[16926] = 8'b1110111;
DRAM[16927] = 8'b1111000;
DRAM[16928] = 8'b1110101;
DRAM[16929] = 8'b1111000;
DRAM[16930] = 8'b1110100;
DRAM[16931] = 8'b1110110;
DRAM[16932] = 8'b1111110;
DRAM[16933] = 8'b1111101;
DRAM[16934] = 8'b1111101;
DRAM[16935] = 8'b10001000;
DRAM[16936] = 8'b10000100;
DRAM[16937] = 8'b10100101;
DRAM[16938] = 8'b11010010;
DRAM[16939] = 8'b11110011;
DRAM[16940] = 8'b11111111;
DRAM[16941] = 8'b11111111;
DRAM[16942] = 8'b11111011;
DRAM[16943] = 8'b11111010;
DRAM[16944] = 8'b11111011;
DRAM[16945] = 8'b11111100;
DRAM[16946] = 8'b11111110;
DRAM[16947] = 8'b11111111;
DRAM[16948] = 8'b11111111;
DRAM[16949] = 8'b11111111;
DRAM[16950] = 8'b11111110;
DRAM[16951] = 8'b11111101;
DRAM[16952] = 8'b11111100;
DRAM[16953] = 8'b11111011;
DRAM[16954] = 8'b11111010;
DRAM[16955] = 8'b11111001;
DRAM[16956] = 8'b11111010;
DRAM[16957] = 8'b11111011;
DRAM[16958] = 8'b11111101;
DRAM[16959] = 8'b11111110;
DRAM[16960] = 8'b11111111;
DRAM[16961] = 8'b11111111;
DRAM[16962] = 8'b11111100;
DRAM[16963] = 8'b11111101;
DRAM[16964] = 8'b11111111;
DRAM[16965] = 8'b11111111;
DRAM[16966] = 8'b11111011;
DRAM[16967] = 8'b11110111;
DRAM[16968] = 8'b11101101;
DRAM[16969] = 8'b11101110;
DRAM[16970] = 8'b11101100;
DRAM[16971] = 8'b11101110;
DRAM[16972] = 8'b11110010;
DRAM[16973] = 8'b11100100;
DRAM[16974] = 8'b10111101;
DRAM[16975] = 8'b10011000;
DRAM[16976] = 8'b1111110;
DRAM[16977] = 8'b1111110;
DRAM[16978] = 8'b1101011;
DRAM[16979] = 8'b1100001;
DRAM[16980] = 8'b1111000;
DRAM[16981] = 8'b10011010;
DRAM[16982] = 8'b10110010;
DRAM[16983] = 8'b11000010;
DRAM[16984] = 8'b11101001;
DRAM[16985] = 8'b11100111;
DRAM[16986] = 8'b11101001;
DRAM[16987] = 8'b11101101;
DRAM[16988] = 8'b11101111;
DRAM[16989] = 8'b11110000;
DRAM[16990] = 8'b11110101;
DRAM[16991] = 8'b11111011;
DRAM[16992] = 8'b11101111;
DRAM[16993] = 8'b11110011;
DRAM[16994] = 8'b11110110;
DRAM[16995] = 8'b11110101;
DRAM[16996] = 8'b11110011;
DRAM[16997] = 8'b11110011;
DRAM[16998] = 8'b11111001;
DRAM[16999] = 8'b11111110;
DRAM[17000] = 8'b11110000;
DRAM[17001] = 8'b11110101;
DRAM[17002] = 8'b11111001;
DRAM[17003] = 8'b11111010;
DRAM[17004] = 8'b11110111;
DRAM[17005] = 8'b11110010;
DRAM[17006] = 8'b11101111;
DRAM[17007] = 8'b11101111;
DRAM[17008] = 8'b11111011;
DRAM[17009] = 8'b11100001;
DRAM[17010] = 8'b11110101;
DRAM[17011] = 8'b11110100;
DRAM[17012] = 8'b11011011;
DRAM[17013] = 8'b11100000;
DRAM[17014] = 8'b11100001;
DRAM[17015] = 8'b11011000;
DRAM[17016] = 8'b11100100;
DRAM[17017] = 8'b11010101;
DRAM[17018] = 8'b11010101;
DRAM[17019] = 8'b11011010;
DRAM[17020] = 8'b11011001;
DRAM[17021] = 8'b11100010;
DRAM[17022] = 8'b11101110;
DRAM[17023] = 8'b11110000;
DRAM[17024] = 8'b11101101;
DRAM[17025] = 8'b11101001;
DRAM[17026] = 8'b11101110;
DRAM[17027] = 8'b11101100;
DRAM[17028] = 8'b11100001;
DRAM[17029] = 8'b11100001;
DRAM[17030] = 8'b11101001;
DRAM[17031] = 8'b11101000;
DRAM[17032] = 8'b11011110;
DRAM[17033] = 8'b11100010;
DRAM[17034] = 8'b11101101;
DRAM[17035] = 8'b11011001;
DRAM[17036] = 8'b11101010;
DRAM[17037] = 8'b11011010;
DRAM[17038] = 8'b11010101;
DRAM[17039] = 8'b11101011;
DRAM[17040] = 8'b11011111;
DRAM[17041] = 8'b11011101;
DRAM[17042] = 8'b11010110;
DRAM[17043] = 8'b11011010;
DRAM[17044] = 8'b11101001;
DRAM[17045] = 8'b11100110;
DRAM[17046] = 8'b11010110;
DRAM[17047] = 8'b11001110;
DRAM[17048] = 8'b11011010;
DRAM[17049] = 8'b11100011;
DRAM[17050] = 8'b11011001;
DRAM[17051] = 8'b11011000;
DRAM[17052] = 8'b11011010;
DRAM[17053] = 8'b11011111;
DRAM[17054] = 8'b11101011;
DRAM[17055] = 8'b11100011;
DRAM[17056] = 8'b11011111;
DRAM[17057] = 8'b11101000;
DRAM[17058] = 8'b11100110;
DRAM[17059] = 8'b11100000;
DRAM[17060] = 8'b11100100;
DRAM[17061] = 8'b11100111;
DRAM[17062] = 8'b11101010;
DRAM[17063] = 8'b11110000;
DRAM[17064] = 8'b11110100;
DRAM[17065] = 8'b11110101;
DRAM[17066] = 8'b11110111;
DRAM[17067] = 8'b11111001;
DRAM[17068] = 8'b11111011;
DRAM[17069] = 8'b11111011;
DRAM[17070] = 8'b11111010;
DRAM[17071] = 8'b11111001;
DRAM[17072] = 8'b11111101;
DRAM[17073] = 8'b11111111;
DRAM[17074] = 8'b11111111;
DRAM[17075] = 8'b11111110;
DRAM[17076] = 8'b11111010;
DRAM[17077] = 8'b11111000;
DRAM[17078] = 8'b11111001;
DRAM[17079] = 8'b11111011;
DRAM[17080] = 8'b11101100;
DRAM[17081] = 8'b11011011;
DRAM[17082] = 8'b11010110;
DRAM[17083] = 8'b10101110;
DRAM[17084] = 8'b1111110;
DRAM[17085] = 8'b1110100;
DRAM[17086] = 8'b1111110;
DRAM[17087] = 8'b10010101;
DRAM[17088] = 8'b10010010;
DRAM[17089] = 8'b10101100;
DRAM[17090] = 8'b11010010;
DRAM[17091] = 8'b11110101;
DRAM[17092] = 8'b11110110;
DRAM[17093] = 8'b11111101;
DRAM[17094] = 8'b11111101;
DRAM[17095] = 8'b11111100;
DRAM[17096] = 8'b11111000;
DRAM[17097] = 8'b11111001;
DRAM[17098] = 8'b11111001;
DRAM[17099] = 8'b11111010;
DRAM[17100] = 8'b11111110;
DRAM[17101] = 8'b11111110;
DRAM[17102] = 8'b11110110;
DRAM[17103] = 8'b11101011;
DRAM[17104] = 8'b11100101;
DRAM[17105] = 8'b11100101;
DRAM[17106] = 8'b11100111;
DRAM[17107] = 8'b11101110;
DRAM[17108] = 8'b11110111;
DRAM[17109] = 8'b11111100;
DRAM[17110] = 8'b11111011;
DRAM[17111] = 8'b11111000;
DRAM[17112] = 8'b11111010;
DRAM[17113] = 8'b11111011;
DRAM[17114] = 8'b11111100;
DRAM[17115] = 8'b11111110;
DRAM[17116] = 8'b11111110;
DRAM[17117] = 8'b11111110;
DRAM[17118] = 8'b11111101;
DRAM[17119] = 8'b11111100;
DRAM[17120] = 8'b11111001;
DRAM[17121] = 8'b11111110;
DRAM[17122] = 8'b11101001;
DRAM[17123] = 8'b10111101;
DRAM[17124] = 8'b10010001;
DRAM[17125] = 8'b1101111;
DRAM[17126] = 8'b1100000;
DRAM[17127] = 8'b1100001;
DRAM[17128] = 8'b1011110;
DRAM[17129] = 8'b1100000;
DRAM[17130] = 8'b1011110;
DRAM[17131] = 8'b1011010;
DRAM[17132] = 8'b1011001;
DRAM[17133] = 8'b1011011;
DRAM[17134] = 8'b1011011;
DRAM[17135] = 8'b1011001;
DRAM[17136] = 8'b1011010;
DRAM[17137] = 8'b1011010;
DRAM[17138] = 8'b1011010;
DRAM[17139] = 8'b1011001;
DRAM[17140] = 8'b1011001;
DRAM[17141] = 8'b1011001;
DRAM[17142] = 8'b1011000;
DRAM[17143] = 8'b1011000;
DRAM[17144] = 8'b1011001;
DRAM[17145] = 8'b1011000;
DRAM[17146] = 8'b1010111;
DRAM[17147] = 8'b1010110;
DRAM[17148] = 8'b1010110;
DRAM[17149] = 8'b1010110;
DRAM[17150] = 8'b1010110;
DRAM[17151] = 8'b1010111;
DRAM[17152] = 8'b1101001;
DRAM[17153] = 8'b1101001;
DRAM[17154] = 8'b1101001;
DRAM[17155] = 8'b1101001;
DRAM[17156] = 8'b1101010;
DRAM[17157] = 8'b1101010;
DRAM[17158] = 8'b1101010;
DRAM[17159] = 8'b1101011;
DRAM[17160] = 8'b1101011;
DRAM[17161] = 8'b1101011;
DRAM[17162] = 8'b1101011;
DRAM[17163] = 8'b1101100;
DRAM[17164] = 8'b1101101;
DRAM[17165] = 8'b1101110;
DRAM[17166] = 8'b1101110;
DRAM[17167] = 8'b1101111;
DRAM[17168] = 8'b1110000;
DRAM[17169] = 8'b1110000;
DRAM[17170] = 8'b1110000;
DRAM[17171] = 8'b1110000;
DRAM[17172] = 8'b1110001;
DRAM[17173] = 8'b1110001;
DRAM[17174] = 8'b1110001;
DRAM[17175] = 8'b1110001;
DRAM[17176] = 8'b1110010;
DRAM[17177] = 8'b1110010;
DRAM[17178] = 8'b1110011;
DRAM[17179] = 8'b1110011;
DRAM[17180] = 8'b1110100;
DRAM[17181] = 8'b1110110;
DRAM[17182] = 8'b1111000;
DRAM[17183] = 8'b1111000;
DRAM[17184] = 8'b1110010;
DRAM[17185] = 8'b1111010;
DRAM[17186] = 8'b1111011;
DRAM[17187] = 8'b1111101;
DRAM[17188] = 8'b10000001;
DRAM[17189] = 8'b10000000;
DRAM[17190] = 8'b10000101;
DRAM[17191] = 8'b10010111;
DRAM[17192] = 8'b10111000;
DRAM[17193] = 8'b11010101;
DRAM[17194] = 8'b11110001;
DRAM[17195] = 8'b11111011;
DRAM[17196] = 8'b11111011;
DRAM[17197] = 8'b11111100;
DRAM[17198] = 8'b11111100;
DRAM[17199] = 8'b11111001;
DRAM[17200] = 8'b11111011;
DRAM[17201] = 8'b11111100;
DRAM[17202] = 8'b11111110;
DRAM[17203] = 8'b11111111;
DRAM[17204] = 8'b11111111;
DRAM[17205] = 8'b11111111;
DRAM[17206] = 8'b11111101;
DRAM[17207] = 8'b11111100;
DRAM[17208] = 8'b11111100;
DRAM[17209] = 8'b11111011;
DRAM[17210] = 8'b11111001;
DRAM[17211] = 8'b11111010;
DRAM[17212] = 8'b11111100;
DRAM[17213] = 8'b11111101;
DRAM[17214] = 8'b11111110;
DRAM[17215] = 8'b11111110;
DRAM[17216] = 8'b11111111;
DRAM[17217] = 8'b11111010;
DRAM[17218] = 8'b11111100;
DRAM[17219] = 8'b11111110;
DRAM[17220] = 8'b11111011;
DRAM[17221] = 8'b11111010;
DRAM[17222] = 8'b11110111;
DRAM[17223] = 8'b11101111;
DRAM[17224] = 8'b11110011;
DRAM[17225] = 8'b11100100;
DRAM[17226] = 8'b11101011;
DRAM[17227] = 8'b11111101;
DRAM[17228] = 8'b11110010;
DRAM[17229] = 8'b11001100;
DRAM[17230] = 8'b10011011;
DRAM[17231] = 8'b1110101;
DRAM[17232] = 8'b10010000;
DRAM[17233] = 8'b1111111;
DRAM[17234] = 8'b1110000;
DRAM[17235] = 8'b1111101;
DRAM[17236] = 8'b10100011;
DRAM[17237] = 8'b11000010;
DRAM[17238] = 8'b11001011;
DRAM[17239] = 8'b11001011;
DRAM[17240] = 8'b11001110;
DRAM[17241] = 8'b11010101;
DRAM[17242] = 8'b11100010;
DRAM[17243] = 8'b11101011;
DRAM[17244] = 8'b11100110;
DRAM[17245] = 8'b11011110;
DRAM[17246] = 8'b11100110;
DRAM[17247] = 8'b11110110;
DRAM[17248] = 8'b11110001;
DRAM[17249] = 8'b11110011;
DRAM[17250] = 8'b11110111;
DRAM[17251] = 8'b11111001;
DRAM[17252] = 8'b11111001;
DRAM[17253] = 8'b11111000;
DRAM[17254] = 8'b11110110;
DRAM[17255] = 8'b11110101;
DRAM[17256] = 8'b11111001;
DRAM[17257] = 8'b11111001;
DRAM[17258] = 8'b11111001;
DRAM[17259] = 8'b11110111;
DRAM[17260] = 8'b11110100;
DRAM[17261] = 8'b11110001;
DRAM[17262] = 8'b11101111;
DRAM[17263] = 8'b11101110;
DRAM[17264] = 8'b11111000;
DRAM[17265] = 8'b11100110;
DRAM[17266] = 8'b11110100;
DRAM[17267] = 8'b11110000;
DRAM[17268] = 8'b11011111;
DRAM[17269] = 8'b11011110;
DRAM[17270] = 8'b11011001;
DRAM[17271] = 8'b11010110;
DRAM[17272] = 8'b11011101;
DRAM[17273] = 8'b11010100;
DRAM[17274] = 8'b11010011;
DRAM[17275] = 8'b11010111;
DRAM[17276] = 8'b11010111;
DRAM[17277] = 8'b11011011;
DRAM[17278] = 8'b11101000;
DRAM[17279] = 8'b11110011;
DRAM[17280] = 8'b11101100;
DRAM[17281] = 8'b11100111;
DRAM[17282] = 8'b11101101;
DRAM[17283] = 8'b11101110;
DRAM[17284] = 8'b11100011;
DRAM[17285] = 8'b11100000;
DRAM[17286] = 8'b11100110;
DRAM[17287] = 8'b11100100;
DRAM[17288] = 8'b11100001;
DRAM[17289] = 8'b11011111;
DRAM[17290] = 8'b11101101;
DRAM[17291] = 8'b11011001;
DRAM[17292] = 8'b11100000;
DRAM[17293] = 8'b11001111;
DRAM[17294] = 8'b11001101;
DRAM[17295] = 8'b11100011;
DRAM[17296] = 8'b11011110;
DRAM[17297] = 8'b11011111;
DRAM[17298] = 8'b11010101;
DRAM[17299] = 8'b11010100;
DRAM[17300] = 8'b11100001;
DRAM[17301] = 8'b11011111;
DRAM[17302] = 8'b11010100;
DRAM[17303] = 8'b11010100;
DRAM[17304] = 8'b11011000;
DRAM[17305] = 8'b11100001;
DRAM[17306] = 8'b11011011;
DRAM[17307] = 8'b11010011;
DRAM[17308] = 8'b11010101;
DRAM[17309] = 8'b11100000;
DRAM[17310] = 8'b11100110;
DRAM[17311] = 8'b11011011;
DRAM[17312] = 8'b11011111;
DRAM[17313] = 8'b11100111;
DRAM[17314] = 8'b11011001;
DRAM[17315] = 8'b11010001;
DRAM[17316] = 8'b11100000;
DRAM[17317] = 8'b11100101;
DRAM[17318] = 8'b11100011;
DRAM[17319] = 8'b11101110;
DRAM[17320] = 8'b11110001;
DRAM[17321] = 8'b11110010;
DRAM[17322] = 8'b11110100;
DRAM[17323] = 8'b11110110;
DRAM[17324] = 8'b11110111;
DRAM[17325] = 8'b11110111;
DRAM[17326] = 8'b11110111;
DRAM[17327] = 8'b11110111;
DRAM[17328] = 8'b11111010;
DRAM[17329] = 8'b11111010;
DRAM[17330] = 8'b11111010;
DRAM[17331] = 8'b11111000;
DRAM[17332] = 8'b11110110;
DRAM[17333] = 8'b11110100;
DRAM[17334] = 8'b11110100;
DRAM[17335] = 8'b11110100;
DRAM[17336] = 8'b11110011;
DRAM[17337] = 8'b11011111;
DRAM[17338] = 8'b11010011;
DRAM[17339] = 8'b10101101;
DRAM[17340] = 8'b10000100;
DRAM[17341] = 8'b1111000;
DRAM[17342] = 8'b10000000;
DRAM[17343] = 8'b10011110;
DRAM[17344] = 8'b10001111;
DRAM[17345] = 8'b10011011;
DRAM[17346] = 8'b10111100;
DRAM[17347] = 8'b11110001;
DRAM[17348] = 8'b11101011;
DRAM[17349] = 8'b11111101;
DRAM[17350] = 8'b11111110;
DRAM[17351] = 8'b11111110;
DRAM[17352] = 8'b11111000;
DRAM[17353] = 8'b11111010;
DRAM[17354] = 8'b11111010;
DRAM[17355] = 8'b11111010;
DRAM[17356] = 8'b11111101;
DRAM[17357] = 8'b11111111;
DRAM[17358] = 8'b11111001;
DRAM[17359] = 8'b11110000;
DRAM[17360] = 8'b11110010;
DRAM[17361] = 8'b11101111;
DRAM[17362] = 8'b11101101;
DRAM[17363] = 8'b11101111;
DRAM[17364] = 8'b11110100;
DRAM[17365] = 8'b11111000;
DRAM[17366] = 8'b11111000;
DRAM[17367] = 8'b11110110;
DRAM[17368] = 8'b11111010;
DRAM[17369] = 8'b11111011;
DRAM[17370] = 8'b11111100;
DRAM[17371] = 8'b11111101;
DRAM[17372] = 8'b11111100;
DRAM[17373] = 8'b11111011;
DRAM[17374] = 8'b11111001;
DRAM[17375] = 8'b11111000;
DRAM[17376] = 8'b11110001;
DRAM[17377] = 8'b11111111;
DRAM[17378] = 8'b11111111;
DRAM[17379] = 8'b11110000;
DRAM[17380] = 8'b11010001;
DRAM[17381] = 8'b10011011;
DRAM[17382] = 8'b1110011;
DRAM[17383] = 8'b1110001;
DRAM[17384] = 8'b1100100;
DRAM[17385] = 8'b1100011;
DRAM[17386] = 8'b1100000;
DRAM[17387] = 8'b1011101;
DRAM[17388] = 8'b1011100;
DRAM[17389] = 8'b1011101;
DRAM[17390] = 8'b1011100;
DRAM[17391] = 8'b1011010;
DRAM[17392] = 8'b1011011;
DRAM[17393] = 8'b1011011;
DRAM[17394] = 8'b1011011;
DRAM[17395] = 8'b1011011;
DRAM[17396] = 8'b1011010;
DRAM[17397] = 8'b1011010;
DRAM[17398] = 8'b1011001;
DRAM[17399] = 8'b1011001;
DRAM[17400] = 8'b1011001;
DRAM[17401] = 8'b1011001;
DRAM[17402] = 8'b1011000;
DRAM[17403] = 8'b1010111;
DRAM[17404] = 8'b1010111;
DRAM[17405] = 8'b1010111;
DRAM[17406] = 8'b1010111;
DRAM[17407] = 8'b1010111;
DRAM[17408] = 8'b1101001;
DRAM[17409] = 8'b1101010;
DRAM[17410] = 8'b1101010;
DRAM[17411] = 8'b1101010;
DRAM[17412] = 8'b1101011;
DRAM[17413] = 8'b1101011;
DRAM[17414] = 8'b1101011;
DRAM[17415] = 8'b1101011;
DRAM[17416] = 8'b1101011;
DRAM[17417] = 8'b1101100;
DRAM[17418] = 8'b1101100;
DRAM[17419] = 8'b1101101;
DRAM[17420] = 8'b1101110;
DRAM[17421] = 8'b1101111;
DRAM[17422] = 8'b1101111;
DRAM[17423] = 8'b1101111;
DRAM[17424] = 8'b1110001;
DRAM[17425] = 8'b1110001;
DRAM[17426] = 8'b1110001;
DRAM[17427] = 8'b1110001;
DRAM[17428] = 8'b1110001;
DRAM[17429] = 8'b1110010;
DRAM[17430] = 8'b1110010;
DRAM[17431] = 8'b1110010;
DRAM[17432] = 8'b1110101;
DRAM[17433] = 8'b1110101;
DRAM[17434] = 8'b1110100;
DRAM[17435] = 8'b1110100;
DRAM[17436] = 8'b1110101;
DRAM[17437] = 8'b1110110;
DRAM[17438] = 8'b1110111;
DRAM[17439] = 8'b1110111;
DRAM[17440] = 8'b1110010;
DRAM[17441] = 8'b1111100;
DRAM[17442] = 8'b1111100;
DRAM[17443] = 8'b1111000;
DRAM[17444] = 8'b1111001;
DRAM[17445] = 8'b1111110;
DRAM[17446] = 8'b10010011;
DRAM[17447] = 8'b10110001;
DRAM[17448] = 8'b11101001;
DRAM[17449] = 8'b11111001;
DRAM[17450] = 8'b11111111;
DRAM[17451] = 8'b11111100;
DRAM[17452] = 8'b11111000;
DRAM[17453] = 8'b11111100;
DRAM[17454] = 8'b11111101;
DRAM[17455] = 8'b11111001;
DRAM[17456] = 8'b11111100;
DRAM[17457] = 8'b11111100;
DRAM[17458] = 8'b11111101;
DRAM[17459] = 8'b11111110;
DRAM[17460] = 8'b11111110;
DRAM[17461] = 8'b11111101;
DRAM[17462] = 8'b11111100;
DRAM[17463] = 8'b11111011;
DRAM[17464] = 8'b11111100;
DRAM[17465] = 8'b11111010;
DRAM[17466] = 8'b11111001;
DRAM[17467] = 8'b11111010;
DRAM[17468] = 8'b11111101;
DRAM[17469] = 8'b11111111;
DRAM[17470] = 8'b11111111;
DRAM[17471] = 8'b11111110;
DRAM[17472] = 8'b11110111;
DRAM[17473] = 8'b11110010;
DRAM[17474] = 8'b11111010;
DRAM[17475] = 8'b11111011;
DRAM[17476] = 8'b11101110;
DRAM[17477] = 8'b11101100;
DRAM[17478] = 8'b11110000;
DRAM[17479] = 8'b11101000;
DRAM[17480] = 8'b11101101;
DRAM[17481] = 8'b11101100;
DRAM[17482] = 8'b11110111;
DRAM[17483] = 8'b11110110;
DRAM[17484] = 8'b11010010;
DRAM[17485] = 8'b10101001;
DRAM[17486] = 8'b10010011;
DRAM[17487] = 8'b10001001;
DRAM[17488] = 8'b10000010;
DRAM[17489] = 8'b1100001;
DRAM[17490] = 8'b1010000;
DRAM[17491] = 8'b1100101;
DRAM[17492] = 8'b10001101;
DRAM[17493] = 8'b10110001;
DRAM[17494] = 8'b11000111;
DRAM[17495] = 8'b11001111;
DRAM[17496] = 8'b11001010;
DRAM[17497] = 8'b11000110;
DRAM[17498] = 8'b11001011;
DRAM[17499] = 8'b11011100;
DRAM[17500] = 8'b11100111;
DRAM[17501] = 8'b11100101;
DRAM[17502] = 8'b11100100;
DRAM[17503] = 8'b11100110;
DRAM[17504] = 8'b11101111;
DRAM[17505] = 8'b11101101;
DRAM[17506] = 8'b11101100;
DRAM[17507] = 8'b11101111;
DRAM[17508] = 8'b11110100;
DRAM[17509] = 8'b11110110;
DRAM[17510] = 8'b11110011;
DRAM[17511] = 8'b11101111;
DRAM[17512] = 8'b11111000;
DRAM[17513] = 8'b11110100;
DRAM[17514] = 8'b11110010;
DRAM[17515] = 8'b11110011;
DRAM[17516] = 8'b11110101;
DRAM[17517] = 8'b11110100;
DRAM[17518] = 8'b11101111;
DRAM[17519] = 8'b11101010;
DRAM[17520] = 8'b11100111;
DRAM[17521] = 8'b11101010;
DRAM[17522] = 8'b11101110;
DRAM[17523] = 8'b11100101;
DRAM[17524] = 8'b11101010;
DRAM[17525] = 8'b11100010;
DRAM[17526] = 8'b11001100;
DRAM[17527] = 8'b11011100;
DRAM[17528] = 8'b11010101;
DRAM[17529] = 8'b11010011;
DRAM[17530] = 8'b11010010;
DRAM[17531] = 8'b11010111;
DRAM[17532] = 8'b11011000;
DRAM[17533] = 8'b11010101;
DRAM[17534] = 8'b11011101;
DRAM[17535] = 8'b11101110;
DRAM[17536] = 8'b11101100;
DRAM[17537] = 8'b11100011;
DRAM[17538] = 8'b11101000;
DRAM[17539] = 8'b11101111;
DRAM[17540] = 8'b11101001;
DRAM[17541] = 8'b11100110;
DRAM[17542] = 8'b11101001;
DRAM[17543] = 8'b11100110;
DRAM[17544] = 8'b11100110;
DRAM[17545] = 8'b11011111;
DRAM[17546] = 8'b11101111;
DRAM[17547] = 8'b11011100;
DRAM[17548] = 8'b11011100;
DRAM[17549] = 8'b11001001;
DRAM[17550] = 8'b11001101;
DRAM[17551] = 8'b11100010;
DRAM[17552] = 8'b11011001;
DRAM[17553] = 8'b11011101;
DRAM[17554] = 8'b11011100;
DRAM[17555] = 8'b11011011;
DRAM[17556] = 8'b11011011;
DRAM[17557] = 8'b11010111;
DRAM[17558] = 8'b11010001;
DRAM[17559] = 8'b11010010;
DRAM[17560] = 8'b11010110;
DRAM[17561] = 8'b11011011;
DRAM[17562] = 8'b11011011;
DRAM[17563] = 8'b11010000;
DRAM[17564] = 8'b11010011;
DRAM[17565] = 8'b11100001;
DRAM[17566] = 8'b11011110;
DRAM[17567] = 8'b11010110;
DRAM[17568] = 8'b11100011;
DRAM[17569] = 8'b11100100;
DRAM[17570] = 8'b11010001;
DRAM[17571] = 8'b11001001;
DRAM[17572] = 8'b11011110;
DRAM[17573] = 8'b11101000;
DRAM[17574] = 8'b11100100;
DRAM[17575] = 8'b11101011;
DRAM[17576] = 8'b11110001;
DRAM[17577] = 8'b11110010;
DRAM[17578] = 8'b11110011;
DRAM[17579] = 8'b11110101;
DRAM[17580] = 8'b11110111;
DRAM[17581] = 8'b11111000;
DRAM[17582] = 8'b11111001;
DRAM[17583] = 8'b11111001;
DRAM[17584] = 8'b11111010;
DRAM[17585] = 8'b11110110;
DRAM[17586] = 8'b11110010;
DRAM[17587] = 8'b11110010;
DRAM[17588] = 8'b11110100;
DRAM[17589] = 8'b11110101;
DRAM[17590] = 8'b11110001;
DRAM[17591] = 8'b11101101;
DRAM[17592] = 8'b11110000;
DRAM[17593] = 8'b11010100;
DRAM[17594] = 8'b11001000;
DRAM[17595] = 8'b10111111;
DRAM[17596] = 8'b10111111;
DRAM[17597] = 8'b10110110;
DRAM[17598] = 8'b10011011;
DRAM[17599] = 8'b10011010;
DRAM[17600] = 8'b10010100;
DRAM[17601] = 8'b10010111;
DRAM[17602] = 8'b10110000;
DRAM[17603] = 8'b11100010;
DRAM[17604] = 8'b11100000;
DRAM[17605] = 8'b11110100;
DRAM[17606] = 8'b11111000;
DRAM[17607] = 8'b11111010;
DRAM[17608] = 8'b11111010;
DRAM[17609] = 8'b11111100;
DRAM[17610] = 8'b11111100;
DRAM[17611] = 8'b11111011;
DRAM[17612] = 8'b11111101;
DRAM[17613] = 8'b11111110;
DRAM[17614] = 8'b11111010;
DRAM[17615] = 8'b11110011;
DRAM[17616] = 8'b11101011;
DRAM[17617] = 8'b11101011;
DRAM[17618] = 8'b11101011;
DRAM[17619] = 8'b11101100;
DRAM[17620] = 8'b11101111;
DRAM[17621] = 8'b11110101;
DRAM[17622] = 8'b11111011;
DRAM[17623] = 8'b11111111;
DRAM[17624] = 8'b11111010;
DRAM[17625] = 8'b11111011;
DRAM[17626] = 8'b11111100;
DRAM[17627] = 8'b11111101;
DRAM[17628] = 8'b11111101;
DRAM[17629] = 8'b11111100;
DRAM[17630] = 8'b11111010;
DRAM[17631] = 8'b11111001;
DRAM[17632] = 8'b11111011;
DRAM[17633] = 8'b11111111;
DRAM[17634] = 8'b11111101;
DRAM[17635] = 8'b11111011;
DRAM[17636] = 8'b11101100;
DRAM[17637] = 8'b10110100;
DRAM[17638] = 8'b10000010;
DRAM[17639] = 8'b1111101;
DRAM[17640] = 8'b1101100;
DRAM[17641] = 8'b1100111;
DRAM[17642] = 8'b1100010;
DRAM[17643] = 8'b1100000;
DRAM[17644] = 8'b1100000;
DRAM[17645] = 8'b1011111;
DRAM[17646] = 8'b1011101;
DRAM[17647] = 8'b1011100;
DRAM[17648] = 8'b1011101;
DRAM[17649] = 8'b1011101;
DRAM[17650] = 8'b1011100;
DRAM[17651] = 8'b1011100;
DRAM[17652] = 8'b1011011;
DRAM[17653] = 8'b1011011;
DRAM[17654] = 8'b1011011;
DRAM[17655] = 8'b1011011;
DRAM[17656] = 8'b1011010;
DRAM[17657] = 8'b1011010;
DRAM[17658] = 8'b1011001;
DRAM[17659] = 8'b1011000;
DRAM[17660] = 8'b1010111;
DRAM[17661] = 8'b1010111;
DRAM[17662] = 8'b1011000;
DRAM[17663] = 8'b1011000;
DRAM[17664] = 8'b1101010;
DRAM[17665] = 8'b1101010;
DRAM[17666] = 8'b1101011;
DRAM[17667] = 8'b1101011;
DRAM[17668] = 8'b1101011;
DRAM[17669] = 8'b1101100;
DRAM[17670] = 8'b1101100;
DRAM[17671] = 8'b1101100;
DRAM[17672] = 8'b1101100;
DRAM[17673] = 8'b1101100;
DRAM[17674] = 8'b1101101;
DRAM[17675] = 8'b1101110;
DRAM[17676] = 8'b1101111;
DRAM[17677] = 8'b1101111;
DRAM[17678] = 8'b1110000;
DRAM[17679] = 8'b1110000;
DRAM[17680] = 8'b1110001;
DRAM[17681] = 8'b1110010;
DRAM[17682] = 8'b1110010;
DRAM[17683] = 8'b1110010;
DRAM[17684] = 8'b1110011;
DRAM[17685] = 8'b1110100;
DRAM[17686] = 8'b1110100;
DRAM[17687] = 8'b1110100;
DRAM[17688] = 8'b1110110;
DRAM[17689] = 8'b1110110;
DRAM[17690] = 8'b1110101;
DRAM[17691] = 8'b1110101;
DRAM[17692] = 8'b1110110;
DRAM[17693] = 8'b1110110;
DRAM[17694] = 8'b1110111;
DRAM[17695] = 8'b1111000;
DRAM[17696] = 8'b1110110;
DRAM[17697] = 8'b1111101;
DRAM[17698] = 8'b1111010;
DRAM[17699] = 8'b1110100;
DRAM[17700] = 8'b1111001;
DRAM[17701] = 8'b10001000;
DRAM[17702] = 8'b10101011;
DRAM[17703] = 8'b11010100;
DRAM[17704] = 8'b11111001;
DRAM[17705] = 8'b11111111;
DRAM[17706] = 8'b11111111;
DRAM[17707] = 8'b11111100;
DRAM[17708] = 8'b11111100;
DRAM[17709] = 8'b11111111;
DRAM[17710] = 8'b11111111;
DRAM[17711] = 8'b11111010;
DRAM[17712] = 8'b11111100;
DRAM[17713] = 8'b11111100;
DRAM[17714] = 8'b11111100;
DRAM[17715] = 8'b11111011;
DRAM[17716] = 8'b11111011;
DRAM[17717] = 8'b11111011;
DRAM[17718] = 8'b11111011;
DRAM[17719] = 8'b11111011;
DRAM[17720] = 8'b11111011;
DRAM[17721] = 8'b11111000;
DRAM[17722] = 8'b11110111;
DRAM[17723] = 8'b11111001;
DRAM[17724] = 8'b11111110;
DRAM[17725] = 8'b11111111;
DRAM[17726] = 8'b11111110;
DRAM[17727] = 8'b11111100;
DRAM[17728] = 8'b11111001;
DRAM[17729] = 8'b11110001;
DRAM[17730] = 8'b11111100;
DRAM[17731] = 8'b11111110;
DRAM[17732] = 8'b11101010;
DRAM[17733] = 8'b11101010;
DRAM[17734] = 8'b11110010;
DRAM[17735] = 8'b11101000;
DRAM[17736] = 8'b11101100;
DRAM[17737] = 8'b11111001;
DRAM[17738] = 8'b11111010;
DRAM[17739] = 8'b11100100;
DRAM[17740] = 8'b11000110;
DRAM[17741] = 8'b10101011;
DRAM[17742] = 8'b10010110;
DRAM[17743] = 8'b10001010;
DRAM[17744] = 8'b10000010;
DRAM[17745] = 8'b1100100;
DRAM[17746] = 8'b1100010;
DRAM[17747] = 8'b1111011;
DRAM[17748] = 8'b10001111;
DRAM[17749] = 8'b10100110;
DRAM[17750] = 8'b11000110;
DRAM[17751] = 8'b11011011;
DRAM[17752] = 8'b11100000;
DRAM[17753] = 8'b11011111;
DRAM[17754] = 8'b11100000;
DRAM[17755] = 8'b11100011;
DRAM[17756] = 8'b11100100;
DRAM[17757] = 8'b11100011;
DRAM[17758] = 8'b11100101;
DRAM[17759] = 8'b11101010;
DRAM[17760] = 8'b11101110;
DRAM[17761] = 8'b11101001;
DRAM[17762] = 8'b11100101;
DRAM[17763] = 8'b11100111;
DRAM[17764] = 8'b11101101;
DRAM[17765] = 8'b11110100;
DRAM[17766] = 8'b11111000;
DRAM[17767] = 8'b11111000;
DRAM[17768] = 8'b11101100;
DRAM[17769] = 8'b11101001;
DRAM[17770] = 8'b11101000;
DRAM[17771] = 8'b11101101;
DRAM[17772] = 8'b11110011;
DRAM[17773] = 8'b11110011;
DRAM[17774] = 8'b11101011;
DRAM[17775] = 8'b11100011;
DRAM[17776] = 8'b11011001;
DRAM[17777] = 8'b11100101;
DRAM[17778] = 8'b11100101;
DRAM[17779] = 8'b11011100;
DRAM[17780] = 8'b11101010;
DRAM[17781] = 8'b11100001;
DRAM[17782] = 8'b11000110;
DRAM[17783] = 8'b11011101;
DRAM[17784] = 8'b11010000;
DRAM[17785] = 8'b11010010;
DRAM[17786] = 8'b11010001;
DRAM[17787] = 8'b11010110;
DRAM[17788] = 8'b11011011;
DRAM[17789] = 8'b11010001;
DRAM[17790] = 8'b11010010;
DRAM[17791] = 8'b11100110;
DRAM[17792] = 8'b11101011;
DRAM[17793] = 8'b11100000;
DRAM[17794] = 8'b11100110;
DRAM[17795] = 8'b11110001;
DRAM[17796] = 8'b11101110;
DRAM[17797] = 8'b11101011;
DRAM[17798] = 8'b11101110;
DRAM[17799] = 8'b11101101;
DRAM[17800] = 8'b11101000;
DRAM[17801] = 8'b11011101;
DRAM[17802] = 8'b11110001;
DRAM[17803] = 8'b11100001;
DRAM[17804] = 8'b11011011;
DRAM[17805] = 8'b11001010;
DRAM[17806] = 8'b11010011;
DRAM[17807] = 8'b11101001;
DRAM[17808] = 8'b11010010;
DRAM[17809] = 8'b11010011;
DRAM[17810] = 8'b11100011;
DRAM[17811] = 8'b11101000;
DRAM[17812] = 8'b11011001;
DRAM[17813] = 8'b11010010;
DRAM[17814] = 8'b11010000;
DRAM[17815] = 8'b11000101;
DRAM[17816] = 8'b11010011;
DRAM[17817] = 8'b11010000;
DRAM[17818] = 8'b11010110;
DRAM[17819] = 8'b11001101;
DRAM[17820] = 8'b11010001;
DRAM[17821] = 8'b11011111;
DRAM[17822] = 8'b11010111;
DRAM[17823] = 8'b11010101;
DRAM[17824] = 8'b11100010;
DRAM[17825] = 8'b11011110;
DRAM[17826] = 8'b11010001;
DRAM[17827] = 8'b11001110;
DRAM[17828] = 8'b11011110;
DRAM[17829] = 8'b11101010;
DRAM[17830] = 8'b11101010;
DRAM[17831] = 8'b11101001;
DRAM[17832] = 8'b11101010;
DRAM[17833] = 8'b11101010;
DRAM[17834] = 8'b11101100;
DRAM[17835] = 8'b11101110;
DRAM[17836] = 8'b11110001;
DRAM[17837] = 8'b11110011;
DRAM[17838] = 8'b11110101;
DRAM[17839] = 8'b11110110;
DRAM[17840] = 8'b11111100;
DRAM[17841] = 8'b11110110;
DRAM[17842] = 8'b11110001;
DRAM[17843] = 8'b11110010;
DRAM[17844] = 8'b11110111;
DRAM[17845] = 8'b11111000;
DRAM[17846] = 8'b11110011;
DRAM[17847] = 8'b11101110;
DRAM[17848] = 8'b11100001;
DRAM[17849] = 8'b11110111;
DRAM[17850] = 8'b11111111;
DRAM[17851] = 8'b11010111;
DRAM[17852] = 8'b10011110;
DRAM[17853] = 8'b1110101;
DRAM[17854] = 8'b1101001;
DRAM[17855] = 8'b10001100;
DRAM[17856] = 8'b10011000;
DRAM[17857] = 8'b10011011;
DRAM[17858] = 8'b10101111;
DRAM[17859] = 8'b11010010;
DRAM[17860] = 8'b11011110;
DRAM[17861] = 8'b11101111;
DRAM[17862] = 8'b11110101;
DRAM[17863] = 8'b11111011;
DRAM[17864] = 8'b11111100;
DRAM[17865] = 8'b11111110;
DRAM[17866] = 8'b11111110;
DRAM[17867] = 8'b11111011;
DRAM[17868] = 8'b11111100;
DRAM[17869] = 8'b11111110;
DRAM[17870] = 8'b11111011;
DRAM[17871] = 8'b11110101;
DRAM[17872] = 8'b11101001;
DRAM[17873] = 8'b11101000;
DRAM[17874] = 8'b11100110;
DRAM[17875] = 8'b11100110;
DRAM[17876] = 8'b11101000;
DRAM[17877] = 8'b11101101;
DRAM[17878] = 8'b11110100;
DRAM[17879] = 8'b11111001;
DRAM[17880] = 8'b11110111;
DRAM[17881] = 8'b11111001;
DRAM[17882] = 8'b11111100;
DRAM[17883] = 8'b11111110;
DRAM[17884] = 8'b11111111;
DRAM[17885] = 8'b11111111;
DRAM[17886] = 8'b11111111;
DRAM[17887] = 8'b11111111;
DRAM[17888] = 8'b11111111;
DRAM[17889] = 8'b11111010;
DRAM[17890] = 8'b11110100;
DRAM[17891] = 8'b11111010;
DRAM[17892] = 8'b11110001;
DRAM[17893] = 8'b11000010;
DRAM[17894] = 8'b10001100;
DRAM[17895] = 8'b1110011;
DRAM[17896] = 8'b1110010;
DRAM[17897] = 8'b1101010;
DRAM[17898] = 8'b1100011;
DRAM[17899] = 8'b1100011;
DRAM[17900] = 8'b1100011;
DRAM[17901] = 8'b1100000;
DRAM[17902] = 8'b1011110;
DRAM[17903] = 8'b1011110;
DRAM[17904] = 8'b1011110;
DRAM[17905] = 8'b1011110;
DRAM[17906] = 8'b1011101;
DRAM[17907] = 8'b1011101;
DRAM[17908] = 8'b1011101;
DRAM[17909] = 8'b1011100;
DRAM[17910] = 8'b1011100;
DRAM[17911] = 8'b1011100;
DRAM[17912] = 8'b1011011;
DRAM[17913] = 8'b1011010;
DRAM[17914] = 8'b1011001;
DRAM[17915] = 8'b1011001;
DRAM[17916] = 8'b1011000;
DRAM[17917] = 8'b1011000;
DRAM[17918] = 8'b1011001;
DRAM[17919] = 8'b1011001;
DRAM[17920] = 8'b1101011;
DRAM[17921] = 8'b1101011;
DRAM[17922] = 8'b1101011;
DRAM[17923] = 8'b1101100;
DRAM[17924] = 8'b1101100;
DRAM[17925] = 8'b1101100;
DRAM[17926] = 8'b1101101;
DRAM[17927] = 8'b1101101;
DRAM[17928] = 8'b1101101;
DRAM[17929] = 8'b1101101;
DRAM[17930] = 8'b1101110;
DRAM[17931] = 8'b1101110;
DRAM[17932] = 8'b1101111;
DRAM[17933] = 8'b1110000;
DRAM[17934] = 8'b1110001;
DRAM[17935] = 8'b1110001;
DRAM[17936] = 8'b1110010;
DRAM[17937] = 8'b1110010;
DRAM[17938] = 8'b1110011;
DRAM[17939] = 8'b1110100;
DRAM[17940] = 8'b1110101;
DRAM[17941] = 8'b1110110;
DRAM[17942] = 8'b1110111;
DRAM[17943] = 8'b1110111;
DRAM[17944] = 8'b1110101;
DRAM[17945] = 8'b1110101;
DRAM[17946] = 8'b1110101;
DRAM[17947] = 8'b1110101;
DRAM[17948] = 8'b1110111;
DRAM[17949] = 8'b1111000;
DRAM[17950] = 8'b1111010;
DRAM[17951] = 8'b1111010;
DRAM[17952] = 8'b1111011;
DRAM[17953] = 8'b10000011;
DRAM[17954] = 8'b10000011;
DRAM[17955] = 8'b10000110;
DRAM[17956] = 8'b10010110;
DRAM[17957] = 8'b10101011;
DRAM[17958] = 8'b11001101;
DRAM[17959] = 8'b11110011;
DRAM[17960] = 8'b11111010;
DRAM[17961] = 8'b11111010;
DRAM[17962] = 8'b11111011;
DRAM[17963] = 8'b11111100;
DRAM[17964] = 8'b11111111;
DRAM[17965] = 8'b11111111;
DRAM[17966] = 8'b11111111;
DRAM[17967] = 8'b11111100;
DRAM[17968] = 8'b11111101;
DRAM[17969] = 8'b11111100;
DRAM[17970] = 8'b11111010;
DRAM[17971] = 8'b11111000;
DRAM[17972] = 8'b11110111;
DRAM[17973] = 8'b11111000;
DRAM[17974] = 8'b11111010;
DRAM[17975] = 8'b11111011;
DRAM[17976] = 8'b11111000;
DRAM[17977] = 8'b11110101;
DRAM[17978] = 8'b11110100;
DRAM[17979] = 8'b11110111;
DRAM[17980] = 8'b11111100;
DRAM[17981] = 8'b11111111;
DRAM[17982] = 8'b11111100;
DRAM[17983] = 8'b11111001;
DRAM[17984] = 8'b11111111;
DRAM[17985] = 8'b11110001;
DRAM[17986] = 8'b11111011;
DRAM[17987] = 8'b11111110;
DRAM[17988] = 8'b11101010;
DRAM[17989] = 8'b11101101;
DRAM[17990] = 8'b11110111;
DRAM[17991] = 8'b11101000;
DRAM[17992] = 8'b11101111;
DRAM[17993] = 8'b11110111;
DRAM[17994] = 8'b11101010;
DRAM[17995] = 8'b11011010;
DRAM[17996] = 8'b11001111;
DRAM[17997] = 8'b10101110;
DRAM[17998] = 8'b10001001;
DRAM[17999] = 8'b10000000;
DRAM[18000] = 8'b1101100;
DRAM[18001] = 8'b1010011;
DRAM[18002] = 8'b1100010;
DRAM[18003] = 8'b10001001;
DRAM[18004] = 8'b10010101;
DRAM[18005] = 8'b10011101;
DRAM[18006] = 8'b10110101;
DRAM[18007] = 8'b11000111;
DRAM[18008] = 8'b11011001;
DRAM[18009] = 8'b11100100;
DRAM[18010] = 8'b11101001;
DRAM[18011] = 8'b11100000;
DRAM[18012] = 8'b11010110;
DRAM[18013] = 8'b11010110;
DRAM[18014] = 8'b11011110;
DRAM[18015] = 8'b11100110;
DRAM[18016] = 8'b11100100;
DRAM[18017] = 8'b11100111;
DRAM[18018] = 8'b11101010;
DRAM[18019] = 8'b11101100;
DRAM[18020] = 8'b11101110;
DRAM[18021] = 8'b11110000;
DRAM[18022] = 8'b11110101;
DRAM[18023] = 8'b11111000;
DRAM[18024] = 8'b11101101;
DRAM[18025] = 8'b11101001;
DRAM[18026] = 8'b11100100;
DRAM[18027] = 8'b11100010;
DRAM[18028] = 8'b11100100;
DRAM[18029] = 8'b11100110;
DRAM[18030] = 8'b11100110;
DRAM[18031] = 8'b11100110;
DRAM[18032] = 8'b11011000;
DRAM[18033] = 8'b11010101;
DRAM[18034] = 8'b11011111;
DRAM[18035] = 8'b11011010;
DRAM[18036] = 8'b11011011;
DRAM[18037] = 8'b11011000;
DRAM[18038] = 8'b11001010;
DRAM[18039] = 8'b11010101;
DRAM[18040] = 8'b11001110;
DRAM[18041] = 8'b11010001;
DRAM[18042] = 8'b11001101;
DRAM[18043] = 8'b11010100;
DRAM[18044] = 8'b11011100;
DRAM[18045] = 8'b11001111;
DRAM[18046] = 8'b11001011;
DRAM[18047] = 8'b11100010;
DRAM[18048] = 8'b11100101;
DRAM[18049] = 8'b11011110;
DRAM[18050] = 8'b11100111;
DRAM[18051] = 8'b11110010;
DRAM[18052] = 8'b11101100;
DRAM[18053] = 8'b11101000;
DRAM[18054] = 8'b11101111;
DRAM[18055] = 8'b11110100;
DRAM[18056] = 8'b11101000;
DRAM[18057] = 8'b11011001;
DRAM[18058] = 8'b11110001;
DRAM[18059] = 8'b11100010;
DRAM[18060] = 8'b11011001;
DRAM[18061] = 8'b11001000;
DRAM[18062] = 8'b11010101;
DRAM[18063] = 8'b11101100;
DRAM[18064] = 8'b11010010;
DRAM[18065] = 8'b11001000;
DRAM[18066] = 8'b11100000;
DRAM[18067] = 8'b11101100;
DRAM[18068] = 8'b11010010;
DRAM[18069] = 8'b11010000;
DRAM[18070] = 8'b11010100;
DRAM[18071] = 8'b10111100;
DRAM[18072] = 8'b11001011;
DRAM[18073] = 8'b11000001;
DRAM[18074] = 8'b11001101;
DRAM[18075] = 8'b11001001;
DRAM[18076] = 8'b11010000;
DRAM[18077] = 8'b11011101;
DRAM[18078] = 8'b11010001;
DRAM[18079] = 8'b11010111;
DRAM[18080] = 8'b11010111;
DRAM[18081] = 8'b11010011;
DRAM[18082] = 8'b11010101;
DRAM[18083] = 8'b11011000;
DRAM[18084] = 8'b11011011;
DRAM[18085] = 8'b11100110;
DRAM[18086] = 8'b11101011;
DRAM[18087] = 8'b11100011;
DRAM[18088] = 8'b11100001;
DRAM[18089] = 8'b11100010;
DRAM[18090] = 8'b11100100;
DRAM[18091] = 8'b11100111;
DRAM[18092] = 8'b11101010;
DRAM[18093] = 8'b11101101;
DRAM[18094] = 8'b11110000;
DRAM[18095] = 8'b11110010;
DRAM[18096] = 8'b11110111;
DRAM[18097] = 8'b11110101;
DRAM[18098] = 8'b11110011;
DRAM[18099] = 8'b11110011;
DRAM[18100] = 8'b11110101;
DRAM[18101] = 8'b11110101;
DRAM[18102] = 8'b11110011;
DRAM[18103] = 8'b11110001;
DRAM[18104] = 8'b11101110;
DRAM[18105] = 8'b11100000;
DRAM[18106] = 8'b11001000;
DRAM[18107] = 8'b10101000;
DRAM[18108] = 8'b10100101;
DRAM[18109] = 8'b10011010;
DRAM[18110] = 8'b1110110;
DRAM[18111] = 8'b1110010;
DRAM[18112] = 8'b10001000;
DRAM[18113] = 8'b10010100;
DRAM[18114] = 8'b10101001;
DRAM[18115] = 8'b10111101;
DRAM[18116] = 8'b11011111;
DRAM[18117] = 8'b11101011;
DRAM[18118] = 8'b11110111;
DRAM[18119] = 8'b11111111;
DRAM[18120] = 8'b11111100;
DRAM[18121] = 8'b11111110;
DRAM[18122] = 8'b11111110;
DRAM[18123] = 8'b11111011;
DRAM[18124] = 8'b11111100;
DRAM[18125] = 8'b11111111;
DRAM[18126] = 8'b11111110;
DRAM[18127] = 8'b11111001;
DRAM[18128] = 8'b11110100;
DRAM[18129] = 8'b11101110;
DRAM[18130] = 8'b11100111;
DRAM[18131] = 8'b11100101;
DRAM[18132] = 8'b11101000;
DRAM[18133] = 8'b11101100;
DRAM[18134] = 8'b11101110;
DRAM[18135] = 8'b11101110;
DRAM[18136] = 8'b11110111;
DRAM[18137] = 8'b11111001;
DRAM[18138] = 8'b11111100;
DRAM[18139] = 8'b11111111;
DRAM[18140] = 8'b11111111;
DRAM[18141] = 8'b11111111;
DRAM[18142] = 8'b11111111;
DRAM[18143] = 8'b11111111;
DRAM[18144] = 8'b11111111;
DRAM[18145] = 8'b11111111;
DRAM[18146] = 8'b11111111;
DRAM[18147] = 8'b11111111;
DRAM[18148] = 8'b11111111;
DRAM[18149] = 8'b11101000;
DRAM[18150] = 8'b10111001;
DRAM[18151] = 8'b10001000;
DRAM[18152] = 8'b1110101;
DRAM[18153] = 8'b1101011;
DRAM[18154] = 8'b1100011;
DRAM[18155] = 8'b1100011;
DRAM[18156] = 8'b1100100;
DRAM[18157] = 8'b1100000;
DRAM[18158] = 8'b1011101;
DRAM[18159] = 8'b1011110;
DRAM[18160] = 8'b1011111;
DRAM[18161] = 8'b1011111;
DRAM[18162] = 8'b1011110;
DRAM[18163] = 8'b1011110;
DRAM[18164] = 8'b1011101;
DRAM[18165] = 8'b1011101;
DRAM[18166] = 8'b1011101;
DRAM[18167] = 8'b1011101;
DRAM[18168] = 8'b1011100;
DRAM[18169] = 8'b1011011;
DRAM[18170] = 8'b1011010;
DRAM[18171] = 8'b1011001;
DRAM[18172] = 8'b1011001;
DRAM[18173] = 8'b1011001;
DRAM[18174] = 8'b1011001;
DRAM[18175] = 8'b1011010;
DRAM[18176] = 8'b1101011;
DRAM[18177] = 8'b1101011;
DRAM[18178] = 8'b1101100;
DRAM[18179] = 8'b1101100;
DRAM[18180] = 8'b1101100;
DRAM[18181] = 8'b1101101;
DRAM[18182] = 8'b1101101;
DRAM[18183] = 8'b1101101;
DRAM[18184] = 8'b1101101;
DRAM[18185] = 8'b1101101;
DRAM[18186] = 8'b1101110;
DRAM[18187] = 8'b1101111;
DRAM[18188] = 8'b1110000;
DRAM[18189] = 8'b1110000;
DRAM[18190] = 8'b1110001;
DRAM[18191] = 8'b1110001;
DRAM[18192] = 8'b1110010;
DRAM[18193] = 8'b1110010;
DRAM[18194] = 8'b1110011;
DRAM[18195] = 8'b1110100;
DRAM[18196] = 8'b1110110;
DRAM[18197] = 8'b1110111;
DRAM[18198] = 8'b1111000;
DRAM[18199] = 8'b1111001;
DRAM[18200] = 8'b1110011;
DRAM[18201] = 8'b1110011;
DRAM[18202] = 8'b1110100;
DRAM[18203] = 8'b1110101;
DRAM[18204] = 8'b1110111;
DRAM[18205] = 8'b1111010;
DRAM[18206] = 8'b1111100;
DRAM[18207] = 8'b1111101;
DRAM[18208] = 8'b1111110;
DRAM[18209] = 8'b10001001;
DRAM[18210] = 8'b10010010;
DRAM[18211] = 8'b10100001;
DRAM[18212] = 8'b10111010;
DRAM[18213] = 8'b11001111;
DRAM[18214] = 8'b11101000;
DRAM[18215] = 8'b11111111;
DRAM[18216] = 8'b11111110;
DRAM[18217] = 8'b11111010;
DRAM[18218] = 8'b11111001;
DRAM[18219] = 8'b11111100;
DRAM[18220] = 8'b11111101;
DRAM[18221] = 8'b11111100;
DRAM[18222] = 8'b11111101;
DRAM[18223] = 8'b11111110;
DRAM[18224] = 8'b11111110;
DRAM[18225] = 8'b11111011;
DRAM[18226] = 8'b11111000;
DRAM[18227] = 8'b11110110;
DRAM[18228] = 8'b11110101;
DRAM[18229] = 8'b11110111;
DRAM[18230] = 8'b11111001;
DRAM[18231] = 8'b11111011;
DRAM[18232] = 8'b11110110;
DRAM[18233] = 8'b11110011;
DRAM[18234] = 8'b11110001;
DRAM[18235] = 8'b11110101;
DRAM[18236] = 8'b11111010;
DRAM[18237] = 8'b11111101;
DRAM[18238] = 8'b11111010;
DRAM[18239] = 8'b11110110;
DRAM[18240] = 8'b11111111;
DRAM[18241] = 8'b11101010;
DRAM[18242] = 8'b11110001;
DRAM[18243] = 8'b11110110;
DRAM[18244] = 8'b11100101;
DRAM[18245] = 8'b11101011;
DRAM[18246] = 8'b11110100;
DRAM[18247] = 8'b11100000;
DRAM[18248] = 8'b11101011;
DRAM[18249] = 8'b11101010;
DRAM[18250] = 8'b11011011;
DRAM[18251] = 8'b11010111;
DRAM[18252] = 8'b11001010;
DRAM[18253] = 8'b10010011;
DRAM[18254] = 8'b1111010;
DRAM[18255] = 8'b10011011;
DRAM[18256] = 8'b1100110;
DRAM[18257] = 8'b1000101;
DRAM[18258] = 8'b1010110;
DRAM[18259] = 8'b10001001;
DRAM[18260] = 8'b10100001;
DRAM[18261] = 8'b10101101;
DRAM[18262] = 8'b11000011;
DRAM[18263] = 8'b11001111;
DRAM[18264] = 8'b11010000;
DRAM[18265] = 8'b11010101;
DRAM[18266] = 8'b11010110;
DRAM[18267] = 8'b11011000;
DRAM[18268] = 8'b11100011;
DRAM[18269] = 8'b11110000;
DRAM[18270] = 8'b11101111;
DRAM[18271] = 8'b11100100;
DRAM[18272] = 8'b11010100;
DRAM[18273] = 8'b11100010;
DRAM[18274] = 8'b11110000;
DRAM[18275] = 8'b11110101;
DRAM[18276] = 8'b11101111;
DRAM[18277] = 8'b11101000;
DRAM[18278] = 8'b11100111;
DRAM[18279] = 8'b11101010;
DRAM[18280] = 8'b11111011;
DRAM[18281] = 8'b11110010;
DRAM[18282] = 8'b11100100;
DRAM[18283] = 8'b11010111;
DRAM[18284] = 8'b11010010;
DRAM[18285] = 8'b11010111;
DRAM[18286] = 8'b11100100;
DRAM[18287] = 8'b11101101;
DRAM[18288] = 8'b11011101;
DRAM[18289] = 8'b11000111;
DRAM[18290] = 8'b11011011;
DRAM[18291] = 8'b11011100;
DRAM[18292] = 8'b11001010;
DRAM[18293] = 8'b11001111;
DRAM[18294] = 8'b11010000;
DRAM[18295] = 8'b11001011;
DRAM[18296] = 8'b11001101;
DRAM[18297] = 8'b11010000;
DRAM[18298] = 8'b11001010;
DRAM[18299] = 8'b11010001;
DRAM[18300] = 8'b11011100;
DRAM[18301] = 8'b11001110;
DRAM[18302] = 8'b11001001;
DRAM[18303] = 8'b11100010;
DRAM[18304] = 8'b11011111;
DRAM[18305] = 8'b11011011;
DRAM[18306] = 8'b11100111;
DRAM[18307] = 8'b11110001;
DRAM[18308] = 8'b11100111;
DRAM[18309] = 8'b11100001;
DRAM[18310] = 8'b11101101;
DRAM[18311] = 8'b11110111;
DRAM[18312] = 8'b11100111;
DRAM[18313] = 8'b11010111;
DRAM[18314] = 8'b11110000;
DRAM[18315] = 8'b11100001;
DRAM[18316] = 8'b11010100;
DRAM[18317] = 8'b11000010;
DRAM[18318] = 8'b11010010;
DRAM[18319] = 8'b11101000;
DRAM[18320] = 8'b11011010;
DRAM[18321] = 8'b11000001;
DRAM[18322] = 8'b11011001;
DRAM[18323] = 8'b11100110;
DRAM[18324] = 8'b11001000;
DRAM[18325] = 8'b11001110;
DRAM[18326] = 8'b11011011;
DRAM[18327] = 8'b10111011;
DRAM[18328] = 8'b11000101;
DRAM[18329] = 8'b10110111;
DRAM[18330] = 8'b11000101;
DRAM[18331] = 8'b11000110;
DRAM[18332] = 8'b11010000;
DRAM[18333] = 8'b11011100;
DRAM[18334] = 8'b11001110;
DRAM[18335] = 8'b11011001;
DRAM[18336] = 8'b11001001;
DRAM[18337] = 8'b11001000;
DRAM[18338] = 8'b11011000;
DRAM[18339] = 8'b11011111;
DRAM[18340] = 8'b11010111;
DRAM[18341] = 8'b11011111;
DRAM[18342] = 8'b11101001;
DRAM[18343] = 8'b11011101;
DRAM[18344] = 8'b11100001;
DRAM[18345] = 8'b11100010;
DRAM[18346] = 8'b11100100;
DRAM[18347] = 8'b11100111;
DRAM[18348] = 8'b11101011;
DRAM[18349] = 8'b11101111;
DRAM[18350] = 8'b11110010;
DRAM[18351] = 8'b11110100;
DRAM[18352] = 8'b11101111;
DRAM[18353] = 8'b11110001;
DRAM[18354] = 8'b11110010;
DRAM[18355] = 8'b11110001;
DRAM[18356] = 8'b11101111;
DRAM[18357] = 8'b11101110;
DRAM[18358] = 8'b11110000;
DRAM[18359] = 8'b11110001;
DRAM[18360] = 8'b11101010;
DRAM[18361] = 8'b11110001;
DRAM[18362] = 8'b11100101;
DRAM[18363] = 8'b10111111;
DRAM[18364] = 8'b10101111;
DRAM[18365] = 8'b10011101;
DRAM[18366] = 8'b1111001;
DRAM[18367] = 8'b1111011;
DRAM[18368] = 8'b1101100;
DRAM[18369] = 8'b10000001;
DRAM[18370] = 8'b10011011;
DRAM[18371] = 8'b10100110;
DRAM[18372] = 8'b11011011;
DRAM[18373] = 8'b11100100;
DRAM[18374] = 8'b11110100;
DRAM[18375] = 8'b11111111;
DRAM[18376] = 8'b11111010;
DRAM[18377] = 8'b11111101;
DRAM[18378] = 8'b11111101;
DRAM[18379] = 8'b11111011;
DRAM[18380] = 8'b11111100;
DRAM[18381] = 8'b11111111;
DRAM[18382] = 8'b11111111;
DRAM[18383] = 8'b11111101;
DRAM[18384] = 8'b11111011;
DRAM[18385] = 8'b11110001;
DRAM[18386] = 8'b11100111;
DRAM[18387] = 8'b11100111;
DRAM[18388] = 8'b11101111;
DRAM[18389] = 8'b11110101;
DRAM[18390] = 8'b11110100;
DRAM[18391] = 8'b11110000;
DRAM[18392] = 8'b11111000;
DRAM[18393] = 8'b11111010;
DRAM[18394] = 8'b11111011;
DRAM[18395] = 8'b11111101;
DRAM[18396] = 8'b11111110;
DRAM[18397] = 8'b11111110;
DRAM[18398] = 8'b11111101;
DRAM[18399] = 8'b11111100;
DRAM[18400] = 8'b11110111;
DRAM[18401] = 8'b11111010;
DRAM[18402] = 8'b11111111;
DRAM[18403] = 8'b11111011;
DRAM[18404] = 8'b11110100;
DRAM[18405] = 8'b11111100;
DRAM[18406] = 8'b11100011;
DRAM[18407] = 8'b10101010;
DRAM[18408] = 8'b1110110;
DRAM[18409] = 8'b1101011;
DRAM[18410] = 8'b1100010;
DRAM[18411] = 8'b1100011;
DRAM[18412] = 8'b1100011;
DRAM[18413] = 8'b1011111;
DRAM[18414] = 8'b1011100;
DRAM[18415] = 8'b1011101;
DRAM[18416] = 8'b1011111;
DRAM[18417] = 8'b1011111;
DRAM[18418] = 8'b1011111;
DRAM[18419] = 8'b1011110;
DRAM[18420] = 8'b1011110;
DRAM[18421] = 8'b1011110;
DRAM[18422] = 8'b1011101;
DRAM[18423] = 8'b1011101;
DRAM[18424] = 8'b1011100;
DRAM[18425] = 8'b1011011;
DRAM[18426] = 8'b1011010;
DRAM[18427] = 8'b1011001;
DRAM[18428] = 8'b1011001;
DRAM[18429] = 8'b1011001;
DRAM[18430] = 8'b1011010;
DRAM[18431] = 8'b1011010;
DRAM[18432] = 8'b1101100;
DRAM[18433] = 8'b1101101;
DRAM[18434] = 8'b1101110;
DRAM[18435] = 8'b1101111;
DRAM[18436] = 8'b1101111;
DRAM[18437] = 8'b1101111;
DRAM[18438] = 8'b1101110;
DRAM[18439] = 8'b1101110;
DRAM[18440] = 8'b1101111;
DRAM[18441] = 8'b1101111;
DRAM[18442] = 8'b1101111;
DRAM[18443] = 8'b1110000;
DRAM[18444] = 8'b1110000;
DRAM[18445] = 8'b1110000;
DRAM[18446] = 8'b1110001;
DRAM[18447] = 8'b1110001;
DRAM[18448] = 8'b1110001;
DRAM[18449] = 8'b1110011;
DRAM[18450] = 8'b1110100;
DRAM[18451] = 8'b1110101;
DRAM[18452] = 8'b1110110;
DRAM[18453] = 8'b1110101;
DRAM[18454] = 8'b1110100;
DRAM[18455] = 8'b1110011;
DRAM[18456] = 8'b1111001;
DRAM[18457] = 8'b1111001;
DRAM[18458] = 8'b1110111;
DRAM[18459] = 8'b1110100;
DRAM[18460] = 8'b1110110;
DRAM[18461] = 8'b1111001;
DRAM[18462] = 8'b1111010;
DRAM[18463] = 8'b1111000;
DRAM[18464] = 8'b10000000;
DRAM[18465] = 8'b10001011;
DRAM[18466] = 8'b10100000;
DRAM[18467] = 8'b10111010;
DRAM[18468] = 8'b11010101;
DRAM[18469] = 8'b11101100;
DRAM[18470] = 8'b11111011;
DRAM[18471] = 8'b11111111;
DRAM[18472] = 8'b11111011;
DRAM[18473] = 8'b11111011;
DRAM[18474] = 8'b11111101;
DRAM[18475] = 8'b11111110;
DRAM[18476] = 8'b11111111;
DRAM[18477] = 8'b11111111;
DRAM[18478] = 8'b11111111;
DRAM[18479] = 8'b11111111;
DRAM[18480] = 8'b11111010;
DRAM[18481] = 8'b11111111;
DRAM[18482] = 8'b11111101;
DRAM[18483] = 8'b11110011;
DRAM[18484] = 8'b11101111;
DRAM[18485] = 8'b11110100;
DRAM[18486] = 8'b11110101;
DRAM[18487] = 8'b11110000;
DRAM[18488] = 8'b11100101;
DRAM[18489] = 8'b11101010;
DRAM[18490] = 8'b11110100;
DRAM[18491] = 8'b11111101;
DRAM[18492] = 8'b11111111;
DRAM[18493] = 8'b11111001;
DRAM[18494] = 8'b11110001;
DRAM[18495] = 8'b11101101;
DRAM[18496] = 8'b11110010;
DRAM[18497] = 8'b11100101;
DRAM[18498] = 8'b11111100;
DRAM[18499] = 8'b11100100;
DRAM[18500] = 8'b11111000;
DRAM[18501] = 8'b11110010;
DRAM[18502] = 8'b11011100;
DRAM[18503] = 8'b11111010;
DRAM[18504] = 8'b11111000;
DRAM[18505] = 8'b11100101;
DRAM[18506] = 8'b11100110;
DRAM[18507] = 8'b11011000;
DRAM[18508] = 8'b10111001;
DRAM[18509] = 8'b10011011;
DRAM[18510] = 8'b10001011;
DRAM[18511] = 8'b10000101;
DRAM[18512] = 8'b1011110;
DRAM[18513] = 8'b1100000;
DRAM[18514] = 8'b10000001;
DRAM[18515] = 8'b10011111;
DRAM[18516] = 8'b10100100;
DRAM[18517] = 8'b10110101;
DRAM[18518] = 8'b11001110;
DRAM[18519] = 8'b11010100;
DRAM[18520] = 8'b11010001;
DRAM[18521] = 8'b11001111;
DRAM[18522] = 8'b11010111;
DRAM[18523] = 8'b11100010;
DRAM[18524] = 8'b11100100;
DRAM[18525] = 8'b11011110;
DRAM[18526] = 8'b11011111;
DRAM[18527] = 8'b11100110;
DRAM[18528] = 8'b11101111;
DRAM[18529] = 8'b11101101;
DRAM[18530] = 8'b11101101;
DRAM[18531] = 8'b11101111;
DRAM[18532] = 8'b11110001;
DRAM[18533] = 8'b11101110;
DRAM[18534] = 8'b11100101;
DRAM[18535] = 8'b11011110;
DRAM[18536] = 8'b11101110;
DRAM[18537] = 8'b11101110;
DRAM[18538] = 8'b11101110;
DRAM[18539] = 8'b11101010;
DRAM[18540] = 8'b11011111;
DRAM[18541] = 8'b11010011;
DRAM[18542] = 8'b11010000;
DRAM[18543] = 8'b11010100;
DRAM[18544] = 8'b11010111;
DRAM[18545] = 8'b11100011;
DRAM[18546] = 8'b10111001;
DRAM[18547] = 8'b11010000;
DRAM[18548] = 8'b11010110;
DRAM[18549] = 8'b11010000;
DRAM[18550] = 8'b11001000;
DRAM[18551] = 8'b11001010;
DRAM[18552] = 8'b11000101;
DRAM[18553] = 8'b11100000;
DRAM[18554] = 8'b11000110;
DRAM[18555] = 8'b11010101;
DRAM[18556] = 8'b11011110;
DRAM[18557] = 8'b10111011;
DRAM[18558] = 8'b11001011;
DRAM[18559] = 8'b11100001;
DRAM[18560] = 8'b11001110;
DRAM[18561] = 8'b11010101;
DRAM[18562] = 8'b11101010;
DRAM[18563] = 8'b11110011;
DRAM[18564] = 8'b11100110;
DRAM[18565] = 8'b11100000;
DRAM[18566] = 8'b11101000;
DRAM[18567] = 8'b11101101;
DRAM[18568] = 8'b11100010;
DRAM[18569] = 8'b11101011;
DRAM[18570] = 8'b11011101;
DRAM[18571] = 8'b11100100;
DRAM[18572] = 8'b11011001;
DRAM[18573] = 8'b11000110;
DRAM[18574] = 8'b11011001;
DRAM[18575] = 8'b11011100;
DRAM[18576] = 8'b11010001;
DRAM[18577] = 8'b11011100;
DRAM[18578] = 8'b11011111;
DRAM[18579] = 8'b11010100;
DRAM[18580] = 8'b11001010;
DRAM[18581] = 8'b11001000;
DRAM[18582] = 8'b11000110;
DRAM[18583] = 8'b11000010;
DRAM[18584] = 8'b11000011;
DRAM[18585] = 8'b10110100;
DRAM[18586] = 8'b11000110;
DRAM[18587] = 8'b11000101;
DRAM[18588] = 8'b11000000;
DRAM[18589] = 8'b11010100;
DRAM[18590] = 8'b11010111;
DRAM[18591] = 8'b11010001;
DRAM[18592] = 8'b11000001;
DRAM[18593] = 8'b10111101;
DRAM[18594] = 8'b11011010;
DRAM[18595] = 8'b11100000;
DRAM[18596] = 8'b11011111;
DRAM[18597] = 8'b11011101;
DRAM[18598] = 8'b11001101;
DRAM[18599] = 8'b11011101;
DRAM[18600] = 8'b11011011;
DRAM[18601] = 8'b11011101;
DRAM[18602] = 8'b11010111;
DRAM[18603] = 8'b11100101;
DRAM[18604] = 8'b11111001;
DRAM[18605] = 8'b11100111;
DRAM[18606] = 8'b11011100;
DRAM[18607] = 8'b11110111;
DRAM[18608] = 8'b11111100;
DRAM[18609] = 8'b11111011;
DRAM[18610] = 8'b11111010;
DRAM[18611] = 8'b11111000;
DRAM[18612] = 8'b11110100;
DRAM[18613] = 8'b11101110;
DRAM[18614] = 8'b11101001;
DRAM[18615] = 8'b11100110;
DRAM[18616] = 8'b11011101;
DRAM[18617] = 8'b11100010;
DRAM[18618] = 8'b11010001;
DRAM[18619] = 8'b11000011;
DRAM[18620] = 8'b10111000;
DRAM[18621] = 8'b10001010;
DRAM[18622] = 8'b1100011;
DRAM[18623] = 8'b1101001;
DRAM[18624] = 8'b1100101;
DRAM[18625] = 8'b10011000;
DRAM[18626] = 8'b10100110;
DRAM[18627] = 8'b10100011;
DRAM[18628] = 8'b10111000;
DRAM[18629] = 8'b11011101;
DRAM[18630] = 8'b11111001;
DRAM[18631] = 8'b11110110;
DRAM[18632] = 8'b11111010;
DRAM[18633] = 8'b11111010;
DRAM[18634] = 8'b11111100;
DRAM[18635] = 8'b11111110;
DRAM[18636] = 8'b11111101;
DRAM[18637] = 8'b11111010;
DRAM[18638] = 8'b11111001;
DRAM[18639] = 8'b11111010;
DRAM[18640] = 8'b11111111;
DRAM[18641] = 8'b11110101;
DRAM[18642] = 8'b11101010;
DRAM[18643] = 8'b11100101;
DRAM[18644] = 8'b11011111;
DRAM[18645] = 8'b11011100;
DRAM[18646] = 8'b11101001;
DRAM[18647] = 8'b11111011;
DRAM[18648] = 8'b11110110;
DRAM[18649] = 8'b11111101;
DRAM[18650] = 8'b11111111;
DRAM[18651] = 8'b11111111;
DRAM[18652] = 8'b11111111;
DRAM[18653] = 8'b11111111;
DRAM[18654] = 8'b11111110;
DRAM[18655] = 8'b11111101;
DRAM[18656] = 8'b11111111;
DRAM[18657] = 8'b11111111;
DRAM[18658] = 8'b11111111;
DRAM[18659] = 8'b11111111;
DRAM[18660] = 8'b11111110;
DRAM[18661] = 8'b11111001;
DRAM[18662] = 8'b11110101;
DRAM[18663] = 8'b11110010;
DRAM[18664] = 8'b10101001;
DRAM[18665] = 8'b10001000;
DRAM[18666] = 8'b1101001;
DRAM[18667] = 8'b1100010;
DRAM[18668] = 8'b1100011;
DRAM[18669] = 8'b1100001;
DRAM[18670] = 8'b1100010;
DRAM[18671] = 8'b1100111;
DRAM[18672] = 8'b1100001;
DRAM[18673] = 8'b1011111;
DRAM[18674] = 8'b1011110;
DRAM[18675] = 8'b1011101;
DRAM[18676] = 8'b1011110;
DRAM[18677] = 8'b1011110;
DRAM[18678] = 8'b1011101;
DRAM[18679] = 8'b1011011;
DRAM[18680] = 8'b1011011;
DRAM[18681] = 8'b1011011;
DRAM[18682] = 8'b1011010;
DRAM[18683] = 8'b1011010;
DRAM[18684] = 8'b1011010;
DRAM[18685] = 8'b1011001;
DRAM[18686] = 8'b1011001;
DRAM[18687] = 8'b1011001;
DRAM[18688] = 8'b1101100;
DRAM[18689] = 8'b1101101;
DRAM[18690] = 8'b1101110;
DRAM[18691] = 8'b1101111;
DRAM[18692] = 8'b1101111;
DRAM[18693] = 8'b1101111;
DRAM[18694] = 8'b1101111;
DRAM[18695] = 8'b1101110;
DRAM[18696] = 8'b1101111;
DRAM[18697] = 8'b1101111;
DRAM[18698] = 8'b1110000;
DRAM[18699] = 8'b1110000;
DRAM[18700] = 8'b1110000;
DRAM[18701] = 8'b1110001;
DRAM[18702] = 8'b1110001;
DRAM[18703] = 8'b1110001;
DRAM[18704] = 8'b1101110;
DRAM[18705] = 8'b1110000;
DRAM[18706] = 8'b1110010;
DRAM[18707] = 8'b1110101;
DRAM[18708] = 8'b1110111;
DRAM[18709] = 8'b1111000;
DRAM[18710] = 8'b1111000;
DRAM[18711] = 8'b1111000;
DRAM[18712] = 8'b1111010;
DRAM[18713] = 8'b1110100;
DRAM[18714] = 8'b1110011;
DRAM[18715] = 8'b1111010;
DRAM[18716] = 8'b10000011;
DRAM[18717] = 8'b10000110;
DRAM[18718] = 8'b10000001;
DRAM[18719] = 8'b1111011;
DRAM[18720] = 8'b1111110;
DRAM[18721] = 8'b10011001;
DRAM[18722] = 8'b11000000;
DRAM[18723] = 8'b11100001;
DRAM[18724] = 8'b11110100;
DRAM[18725] = 8'b11111010;
DRAM[18726] = 8'b11111011;
DRAM[18727] = 8'b11111010;
DRAM[18728] = 8'b11111101;
DRAM[18729] = 8'b11111101;
DRAM[18730] = 8'b11111101;
DRAM[18731] = 8'b11111101;
DRAM[18732] = 8'b11111101;
DRAM[18733] = 8'b11111100;
DRAM[18734] = 8'b11111010;
DRAM[18735] = 8'b11111010;
DRAM[18736] = 8'b11110100;
DRAM[18737] = 8'b11111101;
DRAM[18738] = 8'b11111111;
DRAM[18739] = 8'b11111110;
DRAM[18740] = 8'b11110101;
DRAM[18741] = 8'b11110000;
DRAM[18742] = 8'b11101111;
DRAM[18743] = 8'b11101110;
DRAM[18744] = 8'b11110111;
DRAM[18745] = 8'b11110101;
DRAM[18746] = 8'b11110011;
DRAM[18747] = 8'b11110011;
DRAM[18748] = 8'b11110011;
DRAM[18749] = 8'b11110010;
DRAM[18750] = 8'b11110001;
DRAM[18751] = 8'b11110001;
DRAM[18752] = 8'b11110011;
DRAM[18753] = 8'b11100100;
DRAM[18754] = 8'b11110110;
DRAM[18755] = 8'b11011011;
DRAM[18756] = 8'b11101110;
DRAM[18757] = 8'b11101010;
DRAM[18758] = 8'b11011010;
DRAM[18759] = 8'b11110101;
DRAM[18760] = 8'b11101111;
DRAM[18761] = 8'b11100010;
DRAM[18762] = 8'b11001010;
DRAM[18763] = 8'b11001100;
DRAM[18764] = 8'b10111010;
DRAM[18765] = 8'b10000101;
DRAM[18766] = 8'b10100011;
DRAM[18767] = 8'b1111011;
DRAM[18768] = 8'b1101100;
DRAM[18769] = 8'b1100010;
DRAM[18770] = 8'b1110100;
DRAM[18771] = 8'b10001101;
DRAM[18772] = 8'b10011001;
DRAM[18773] = 8'b10101100;
DRAM[18774] = 8'b10111101;
DRAM[18775] = 8'b10111011;
DRAM[18776] = 8'b11010101;
DRAM[18777] = 8'b11001100;
DRAM[18778] = 8'b11001001;
DRAM[18779] = 8'b11010110;
DRAM[18780] = 8'b11100110;
DRAM[18781] = 8'b11101101;
DRAM[18782] = 8'b11101010;
DRAM[18783] = 8'b11100110;
DRAM[18784] = 8'b11011111;
DRAM[18785] = 8'b11011111;
DRAM[18786] = 8'b11100000;
DRAM[18787] = 8'b11100100;
DRAM[18788] = 8'b11101000;
DRAM[18789] = 8'b11101011;
DRAM[18790] = 8'b11101010;
DRAM[18791] = 8'b11101000;
DRAM[18792] = 8'b11011100;
DRAM[18793] = 8'b11011111;
DRAM[18794] = 8'b11101000;
DRAM[18795] = 8'b11101111;
DRAM[18796] = 8'b11101100;
DRAM[18797] = 8'b11011110;
DRAM[18798] = 8'b11010011;
DRAM[18799] = 8'b11001111;
DRAM[18800] = 8'b11010001;
DRAM[18801] = 8'b11010100;
DRAM[18802] = 8'b11000001;
DRAM[18803] = 8'b11000000;
DRAM[18804] = 8'b11010011;
DRAM[18805] = 8'b11001101;
DRAM[18806] = 8'b11010000;
DRAM[18807] = 8'b11010101;
DRAM[18808] = 8'b11001101;
DRAM[18809] = 8'b11011101;
DRAM[18810] = 8'b11001010;
DRAM[18811] = 8'b11001110;
DRAM[18812] = 8'b11011010;
DRAM[18813] = 8'b11000110;
DRAM[18814] = 8'b11000101;
DRAM[18815] = 8'b11010110;
DRAM[18816] = 8'b11010010;
DRAM[18817] = 8'b11010100;
DRAM[18818] = 8'b11100011;
DRAM[18819] = 8'b11101011;
DRAM[18820] = 8'b11100001;
DRAM[18821] = 8'b11011110;
DRAM[18822] = 8'b11100111;
DRAM[18823] = 8'b11101010;
DRAM[18824] = 8'b11100001;
DRAM[18825] = 8'b11101001;
DRAM[18826] = 8'b11011110;
DRAM[18827] = 8'b11100011;
DRAM[18828] = 8'b11011001;
DRAM[18829] = 8'b11001010;
DRAM[18830] = 8'b11011011;
DRAM[18831] = 8'b11011110;
DRAM[18832] = 8'b11010011;
DRAM[18833] = 8'b11011011;
DRAM[18834] = 8'b11011001;
DRAM[18835] = 8'b11001100;
DRAM[18836] = 8'b11000011;
DRAM[18837] = 8'b11000100;
DRAM[18838] = 8'b11000101;
DRAM[18839] = 8'b11000010;
DRAM[18840] = 8'b11000000;
DRAM[18841] = 8'b10101101;
DRAM[18842] = 8'b10111011;
DRAM[18843] = 8'b11000100;
DRAM[18844] = 8'b11001101;
DRAM[18845] = 8'b11011111;
DRAM[18846] = 8'b11010001;
DRAM[18847] = 8'b10111100;
DRAM[18848] = 8'b10111110;
DRAM[18849] = 8'b11001111;
DRAM[18850] = 8'b11100101;
DRAM[18851] = 8'b11010000;
DRAM[18852] = 8'b11001011;
DRAM[18853] = 8'b11011101;
DRAM[18854] = 8'b11010001;
DRAM[18855] = 8'b11001101;
DRAM[18856] = 8'b11011100;
DRAM[18857] = 8'b11001110;
DRAM[18858] = 8'b11010010;
DRAM[18859] = 8'b11100110;
DRAM[18860] = 8'b11101101;
DRAM[18861] = 8'b11101011;
DRAM[18862] = 8'b11101010;
DRAM[18863] = 8'b11101011;
DRAM[18864] = 8'b11101011;
DRAM[18865] = 8'b11101101;
DRAM[18866] = 8'b11110001;
DRAM[18867] = 8'b11110100;
DRAM[18868] = 8'b11110110;
DRAM[18869] = 8'b11110101;
DRAM[18870] = 8'b11110011;
DRAM[18871] = 8'b11110010;
DRAM[18872] = 8'b11101000;
DRAM[18873] = 8'b11010111;
DRAM[18874] = 8'b11001111;
DRAM[18875] = 8'b11000111;
DRAM[18876] = 8'b10110001;
DRAM[18877] = 8'b10100001;
DRAM[18878] = 8'b10011001;
DRAM[18879] = 8'b10001110;
DRAM[18880] = 8'b1101001;
DRAM[18881] = 8'b10000110;
DRAM[18882] = 8'b10011111;
DRAM[18883] = 8'b10100101;
DRAM[18884] = 8'b10101110;
DRAM[18885] = 8'b11000101;
DRAM[18886] = 8'b11100011;
DRAM[18887] = 8'b11111111;
DRAM[18888] = 8'b11111100;
DRAM[18889] = 8'b11111001;
DRAM[18890] = 8'b11110111;
DRAM[18891] = 8'b11111010;
DRAM[18892] = 8'b11111101;
DRAM[18893] = 8'b11111101;
DRAM[18894] = 8'b11111011;
DRAM[18895] = 8'b11111001;
DRAM[18896] = 8'b11111111;
DRAM[18897] = 8'b11111001;
DRAM[18898] = 8'b11110101;
DRAM[18899] = 8'b11110011;
DRAM[18900] = 8'b11101010;
DRAM[18901] = 8'b11011101;
DRAM[18902] = 8'b11011101;
DRAM[18903] = 8'b11100111;
DRAM[18904] = 8'b11111000;
DRAM[18905] = 8'b11110111;
DRAM[18906] = 8'b11110101;
DRAM[18907] = 8'b11111000;
DRAM[18908] = 8'b11111110;
DRAM[18909] = 8'b11111111;
DRAM[18910] = 8'b11111111;
DRAM[18911] = 8'b11111100;
DRAM[18912] = 8'b11111101;
DRAM[18913] = 8'b11111110;
DRAM[18914] = 8'b11111111;
DRAM[18915] = 8'b11111111;
DRAM[18916] = 8'b11111110;
DRAM[18917] = 8'b11111100;
DRAM[18918] = 8'b11111000;
DRAM[18919] = 8'b11110110;
DRAM[18920] = 8'b11010110;
DRAM[18921] = 8'b10110000;
DRAM[18922] = 8'b10000110;
DRAM[18923] = 8'b1110010;
DRAM[18924] = 8'b1110000;
DRAM[18925] = 8'b1101101;
DRAM[18926] = 8'b1100110;
DRAM[18927] = 8'b1100000;
DRAM[18928] = 8'b1011111;
DRAM[18929] = 8'b1011110;
DRAM[18930] = 8'b1011100;
DRAM[18931] = 8'b1011100;
DRAM[18932] = 8'b1011101;
DRAM[18933] = 8'b1011110;
DRAM[18934] = 8'b1011101;
DRAM[18935] = 8'b1011011;
DRAM[18936] = 8'b1011011;
DRAM[18937] = 8'b1011011;
DRAM[18938] = 8'b1011011;
DRAM[18939] = 8'b1011010;
DRAM[18940] = 8'b1011010;
DRAM[18941] = 8'b1011010;
DRAM[18942] = 8'b1011001;
DRAM[18943] = 8'b1011001;
DRAM[18944] = 8'b1101101;
DRAM[18945] = 8'b1101110;
DRAM[18946] = 8'b1101111;
DRAM[18947] = 8'b1101111;
DRAM[18948] = 8'b1110000;
DRAM[18949] = 8'b1110000;
DRAM[18950] = 8'b1101111;
DRAM[18951] = 8'b1101111;
DRAM[18952] = 8'b1110000;
DRAM[18953] = 8'b1110000;
DRAM[18954] = 8'b1110000;
DRAM[18955] = 8'b1110001;
DRAM[18956] = 8'b1110001;
DRAM[18957] = 8'b1110001;
DRAM[18958] = 8'b1110010;
DRAM[18959] = 8'b1110010;
DRAM[18960] = 8'b1101111;
DRAM[18961] = 8'b1110000;
DRAM[18962] = 8'b1110011;
DRAM[18963] = 8'b1110101;
DRAM[18964] = 8'b1110111;
DRAM[18965] = 8'b1111001;
DRAM[18966] = 8'b1111001;
DRAM[18967] = 8'b1111010;
DRAM[18968] = 8'b1111100;
DRAM[18969] = 8'b1110111;
DRAM[18970] = 8'b1111000;
DRAM[18971] = 8'b1111111;
DRAM[18972] = 8'b10000001;
DRAM[18973] = 8'b1111101;
DRAM[18974] = 8'b1111110;
DRAM[18975] = 8'b10000011;
DRAM[18976] = 8'b10011111;
DRAM[18977] = 8'b10111110;
DRAM[18978] = 8'b11100111;
DRAM[18979] = 8'b11111111;
DRAM[18980] = 8'b11111111;
DRAM[18981] = 8'b11111111;
DRAM[18982] = 8'b11111010;
DRAM[18983] = 8'b11111000;
DRAM[18984] = 8'b11111110;
DRAM[18985] = 8'b11111110;
DRAM[18986] = 8'b11111110;
DRAM[18987] = 8'b11111110;
DRAM[18988] = 8'b11111101;
DRAM[18989] = 8'b11111100;
DRAM[18990] = 8'b11111010;
DRAM[18991] = 8'b11111001;
DRAM[18992] = 8'b11111011;
DRAM[18993] = 8'b11110101;
DRAM[18994] = 8'b11101111;
DRAM[18995] = 8'b11101101;
DRAM[18996] = 8'b11101011;
DRAM[18997] = 8'b11101010;
DRAM[18998] = 8'b11101101;
DRAM[18999] = 8'b11110011;
DRAM[19000] = 8'b11111001;
DRAM[19001] = 8'b11110110;
DRAM[19002] = 8'b11110010;
DRAM[19003] = 8'b11110001;
DRAM[19004] = 8'b11110100;
DRAM[19005] = 8'b11111000;
DRAM[19006] = 8'b11111011;
DRAM[19007] = 8'b11111100;
DRAM[19008] = 8'b11101010;
DRAM[19009] = 8'b11100001;
DRAM[19010] = 8'b11110110;
DRAM[19011] = 8'b11011111;
DRAM[19012] = 8'b11101101;
DRAM[19013] = 8'b11101010;
DRAM[19014] = 8'b11011111;
DRAM[19015] = 8'b11110011;
DRAM[19016] = 8'b11101010;
DRAM[19017] = 8'b11011111;
DRAM[19018] = 8'b10101000;
DRAM[19019] = 8'b11011000;
DRAM[19020] = 8'b10010010;
DRAM[19021] = 8'b10010111;
DRAM[19022] = 8'b10010101;
DRAM[19023] = 8'b1110110;
DRAM[19024] = 8'b1000010;
DRAM[19025] = 8'b1010001;
DRAM[19026] = 8'b1110011;
DRAM[19027] = 8'b10001010;
DRAM[19028] = 8'b10001111;
DRAM[19029] = 8'b10100101;
DRAM[19030] = 8'b11001011;
DRAM[19031] = 8'b11100011;
DRAM[19032] = 8'b11010111;
DRAM[19033] = 8'b11011100;
DRAM[19034] = 8'b11011110;
DRAM[19035] = 8'b11011100;
DRAM[19036] = 8'b11011100;
DRAM[19037] = 8'b11100011;
DRAM[19038] = 8'b11101010;
DRAM[19039] = 8'b11101101;
DRAM[19040] = 8'b11100110;
DRAM[19041] = 8'b11100110;
DRAM[19042] = 8'b11100110;
DRAM[19043] = 8'b11100101;
DRAM[19044] = 8'b11100101;
DRAM[19045] = 8'b11100110;
DRAM[19046] = 8'b11101000;
DRAM[19047] = 8'b11101011;
DRAM[19048] = 8'b11101000;
DRAM[19049] = 8'b11100010;
DRAM[19050] = 8'b11100000;
DRAM[19051] = 8'b11100100;
DRAM[19052] = 8'b11100101;
DRAM[19053] = 8'b11011111;
DRAM[19054] = 8'b11011000;
DRAM[19055] = 8'b11010100;
DRAM[19056] = 8'b11001110;
DRAM[19057] = 8'b11001001;
DRAM[19058] = 8'b11001110;
DRAM[19059] = 8'b10110011;
DRAM[19060] = 8'b11001001;
DRAM[19061] = 8'b11000111;
DRAM[19062] = 8'b11010000;
DRAM[19063] = 8'b11011010;
DRAM[19064] = 8'b11001011;
DRAM[19065] = 8'b11001110;
DRAM[19066] = 8'b11000111;
DRAM[19067] = 8'b10111101;
DRAM[19068] = 8'b11001011;
DRAM[19069] = 8'b11001010;
DRAM[19070] = 8'b10110110;
DRAM[19071] = 8'b11000001;
DRAM[19072] = 8'b11010101;
DRAM[19073] = 8'b11010000;
DRAM[19074] = 8'b11011000;
DRAM[19075] = 8'b11100000;
DRAM[19076] = 8'b11011011;
DRAM[19077] = 8'b11011100;
DRAM[19078] = 8'b11100100;
DRAM[19079] = 8'b11100101;
DRAM[19080] = 8'b11011101;
DRAM[19081] = 8'b11100011;
DRAM[19082] = 8'b11011100;
DRAM[19083] = 8'b11011111;
DRAM[19084] = 8'b11010110;
DRAM[19085] = 8'b11001100;
DRAM[19086] = 8'b11011000;
DRAM[19087] = 8'b11011100;
DRAM[19088] = 8'b11010101;
DRAM[19089] = 8'b11011000;
DRAM[19090] = 8'b11010001;
DRAM[19091] = 8'b11000011;
DRAM[19092] = 8'b10111100;
DRAM[19093] = 8'b11000010;
DRAM[19094] = 8'b11001001;
DRAM[19095] = 8'b11001001;
DRAM[19096] = 8'b10101100;
DRAM[19097] = 8'b10101010;
DRAM[19098] = 8'b11000001;
DRAM[19099] = 8'b11000100;
DRAM[19100] = 8'b11000011;
DRAM[19101] = 8'b11001100;
DRAM[19102] = 8'b11000010;
DRAM[19103] = 8'b10111001;
DRAM[19104] = 8'b11001000;
DRAM[19105] = 8'b11000101;
DRAM[19106] = 8'b11010000;
DRAM[19107] = 8'b11001100;
DRAM[19108] = 8'b11000101;
DRAM[19109] = 8'b11000101;
DRAM[19110] = 8'b11000010;
DRAM[19111] = 8'b11010000;
DRAM[19112] = 8'b11100000;
DRAM[19113] = 8'b11001110;
DRAM[19114] = 8'b11011101;
DRAM[19115] = 8'b11101001;
DRAM[19116] = 8'b11011001;
DRAM[19117] = 8'b11011110;
DRAM[19118] = 8'b11101011;
DRAM[19119] = 8'b11011101;
DRAM[19120] = 8'b11101000;
DRAM[19121] = 8'b11101011;
DRAM[19122] = 8'b11110000;
DRAM[19123] = 8'b11110011;
DRAM[19124] = 8'b11110100;
DRAM[19125] = 8'b11110010;
DRAM[19126] = 8'b11101111;
DRAM[19127] = 8'b11101100;
DRAM[19128] = 8'b11011101;
DRAM[19129] = 8'b11100011;
DRAM[19130] = 8'b11001101;
DRAM[19131] = 8'b10110101;
DRAM[19132] = 8'b10101111;
DRAM[19133] = 8'b10010110;
DRAM[19134] = 8'b1110011;
DRAM[19135] = 8'b1101011;
DRAM[19136] = 8'b1110111;
DRAM[19137] = 8'b1110111;
DRAM[19138] = 8'b10010101;
DRAM[19139] = 8'b10011100;
DRAM[19140] = 8'b10101111;
DRAM[19141] = 8'b11010001;
DRAM[19142] = 8'b11011101;
DRAM[19143] = 8'b11111101;
DRAM[19144] = 8'b11111110;
DRAM[19145] = 8'b11111000;
DRAM[19146] = 8'b11110100;
DRAM[19147] = 8'b11110101;
DRAM[19148] = 8'b11111011;
DRAM[19149] = 8'b11111111;
DRAM[19150] = 8'b11111101;
DRAM[19151] = 8'b11111000;
DRAM[19152] = 8'b11111010;
DRAM[19153] = 8'b11110111;
DRAM[19154] = 8'b11111000;
DRAM[19155] = 8'b11111001;
DRAM[19156] = 8'b11101111;
DRAM[19157] = 8'b11011111;
DRAM[19158] = 8'b11011001;
DRAM[19159] = 8'b11011100;
DRAM[19160] = 8'b11101110;
DRAM[19161] = 8'b11101110;
DRAM[19162] = 8'b11110001;
DRAM[19163] = 8'b11110111;
DRAM[19164] = 8'b11111100;
DRAM[19165] = 8'b11111110;
DRAM[19166] = 8'b11111110;
DRAM[19167] = 8'b11111101;
DRAM[19168] = 8'b11111011;
DRAM[19169] = 8'b11111100;
DRAM[19170] = 8'b11111110;
DRAM[19171] = 8'b11111111;
DRAM[19172] = 8'b11111111;
DRAM[19173] = 8'b11111110;
DRAM[19174] = 8'b11111100;
DRAM[19175] = 8'b11111011;
DRAM[19176] = 8'b11111111;
DRAM[19177] = 8'b11010110;
DRAM[19178] = 8'b10011011;
DRAM[19179] = 8'b1110001;
DRAM[19180] = 8'b1100110;
DRAM[19181] = 8'b1101001;
DRAM[19182] = 8'b1100110;
DRAM[19183] = 8'b1011101;
DRAM[19184] = 8'b1100000;
DRAM[19185] = 8'b1011110;
DRAM[19186] = 8'b1011100;
DRAM[19187] = 8'b1011100;
DRAM[19188] = 8'b1011101;
DRAM[19189] = 8'b1011110;
DRAM[19190] = 8'b1011101;
DRAM[19191] = 8'b1011100;
DRAM[19192] = 8'b1011100;
DRAM[19193] = 8'b1011100;
DRAM[19194] = 8'b1011011;
DRAM[19195] = 8'b1011011;
DRAM[19196] = 8'b1011011;
DRAM[19197] = 8'b1011010;
DRAM[19198] = 8'b1011010;
DRAM[19199] = 8'b1011010;
DRAM[19200] = 8'b1101110;
DRAM[19201] = 8'b1101110;
DRAM[19202] = 8'b1101111;
DRAM[19203] = 8'b1110000;
DRAM[19204] = 8'b1110001;
DRAM[19205] = 8'b1110001;
DRAM[19206] = 8'b1110000;
DRAM[19207] = 8'b1110000;
DRAM[19208] = 8'b1110001;
DRAM[19209] = 8'b1110001;
DRAM[19210] = 8'b1110001;
DRAM[19211] = 8'b1110001;
DRAM[19212] = 8'b1110010;
DRAM[19213] = 8'b1110010;
DRAM[19214] = 8'b1110010;
DRAM[19215] = 8'b1110011;
DRAM[19216] = 8'b1110100;
DRAM[19217] = 8'b1110101;
DRAM[19218] = 8'b1110101;
DRAM[19219] = 8'b1110110;
DRAM[19220] = 8'b1110111;
DRAM[19221] = 8'b1111000;
DRAM[19222] = 8'b1111000;
DRAM[19223] = 8'b1111000;
DRAM[19224] = 8'b1111000;
DRAM[19225] = 8'b1111010;
DRAM[19226] = 8'b10000000;
DRAM[19227] = 8'b10000000;
DRAM[19228] = 8'b1110111;
DRAM[19229] = 8'b1110111;
DRAM[19230] = 8'b10010000;
DRAM[19231] = 8'b10101111;
DRAM[19232] = 8'b11011011;
DRAM[19233] = 8'b11101011;
DRAM[19234] = 8'b11111101;
DRAM[19235] = 8'b11111111;
DRAM[19236] = 8'b11111110;
DRAM[19237] = 8'b11111001;
DRAM[19238] = 8'b11111010;
DRAM[19239] = 8'b11111110;
DRAM[19240] = 8'b11111101;
DRAM[19241] = 8'b11111110;
DRAM[19242] = 8'b11111111;
DRAM[19243] = 8'b11111111;
DRAM[19244] = 8'b11111111;
DRAM[19245] = 8'b11111111;
DRAM[19246] = 8'b11111111;
DRAM[19247] = 8'b11111110;
DRAM[19248] = 8'b11111111;
DRAM[19249] = 8'b11101011;
DRAM[19250] = 8'b11011110;
DRAM[19251] = 8'b11100100;
DRAM[19252] = 8'b11101111;
DRAM[19253] = 8'b11110000;
DRAM[19254] = 8'b11101110;
DRAM[19255] = 8'b11101110;
DRAM[19256] = 8'b11101110;
DRAM[19257] = 8'b11110010;
DRAM[19258] = 8'b11110101;
DRAM[19259] = 8'b11111000;
DRAM[19260] = 8'b11111100;
DRAM[19261] = 8'b11111110;
DRAM[19262] = 8'b11111001;
DRAM[19263] = 8'b11110010;
DRAM[19264] = 8'b11010011;
DRAM[19265] = 8'b11011000;
DRAM[19266] = 8'b11110111;
DRAM[19267] = 8'b11100111;
DRAM[19268] = 8'b11101110;
DRAM[19269] = 8'b11100111;
DRAM[19270] = 8'b11100100;
DRAM[19271] = 8'b11101101;
DRAM[19272] = 8'b11110010;
DRAM[19273] = 8'b11001011;
DRAM[19274] = 8'b10110100;
DRAM[19275] = 8'b11010110;
DRAM[19276] = 8'b1111010;
DRAM[19277] = 8'b10101010;
DRAM[19278] = 8'b1111001;
DRAM[19279] = 8'b1110000;
DRAM[19280] = 8'b1100110;
DRAM[19281] = 8'b1100101;
DRAM[19282] = 8'b1110001;
DRAM[19283] = 8'b10001010;
DRAM[19284] = 8'b10100101;
DRAM[19285] = 8'b10111011;
DRAM[19286] = 8'b11000110;
DRAM[19287] = 8'b11000101;
DRAM[19288] = 8'b11010100;
DRAM[19289] = 8'b11100011;
DRAM[19290] = 8'b11101000;
DRAM[19291] = 8'b11011101;
DRAM[19292] = 8'b11010100;
DRAM[19293] = 8'b11011001;
DRAM[19294] = 8'b11100100;
DRAM[19295] = 8'b11101001;
DRAM[19296] = 8'b11110000;
DRAM[19297] = 8'b11110010;
DRAM[19298] = 8'b11110010;
DRAM[19299] = 8'b11101101;
DRAM[19300] = 8'b11100110;
DRAM[19301] = 8'b11100011;
DRAM[19302] = 8'b11100101;
DRAM[19303] = 8'b11101000;
DRAM[19304] = 8'b11101111;
DRAM[19305] = 8'b11100001;
DRAM[19306] = 8'b11010110;
DRAM[19307] = 8'b11011000;
DRAM[19308] = 8'b11011111;
DRAM[19309] = 8'b11100001;
DRAM[19310] = 8'b11011111;
DRAM[19311] = 8'b11011110;
DRAM[19312] = 8'b11010001;
DRAM[19313] = 8'b11001001;
DRAM[19314] = 8'b11010111;
DRAM[19315] = 8'b10110111;
DRAM[19316] = 8'b10111011;
DRAM[19317] = 8'b11000011;
DRAM[19318] = 8'b11000100;
DRAM[19319] = 8'b11010011;
DRAM[19320] = 8'b11000110;
DRAM[19321] = 8'b10111111;
DRAM[19322] = 8'b11001001;
DRAM[19323] = 8'b10110000;
DRAM[19324] = 8'b10111011;
DRAM[19325] = 8'b11001011;
DRAM[19326] = 8'b10101100;
DRAM[19327] = 8'b10110111;
DRAM[19328] = 8'b11010100;
DRAM[19329] = 8'b11001011;
DRAM[19330] = 8'b11010000;
DRAM[19331] = 8'b11011001;
DRAM[19332] = 8'b11010111;
DRAM[19333] = 8'b11011010;
DRAM[19334] = 8'b11100000;
DRAM[19335] = 8'b11011101;
DRAM[19336] = 8'b11011000;
DRAM[19337] = 8'b11011100;
DRAM[19338] = 8'b11011010;
DRAM[19339] = 8'b11011000;
DRAM[19340] = 8'b11010000;
DRAM[19341] = 8'b11001011;
DRAM[19342] = 8'b11010001;
DRAM[19343] = 8'b11010101;
DRAM[19344] = 8'b11010111;
DRAM[19345] = 8'b11010110;
DRAM[19346] = 8'b11001011;
DRAM[19347] = 8'b10111100;
DRAM[19348] = 8'b10111001;
DRAM[19349] = 8'b11000100;
DRAM[19350] = 8'b11001110;
DRAM[19351] = 8'b11001111;
DRAM[19352] = 8'b10101010;
DRAM[19353] = 8'b10110000;
DRAM[19354] = 8'b11000110;
DRAM[19355] = 8'b11000000;
DRAM[19356] = 8'b10111000;
DRAM[19357] = 8'b10111101;
DRAM[19358] = 8'b10111000;
DRAM[19359] = 8'b10111101;
DRAM[19360] = 8'b11001110;
DRAM[19361] = 8'b10111011;
DRAM[19362] = 8'b10111011;
DRAM[19363] = 8'b11000101;
DRAM[19364] = 8'b11000110;
DRAM[19365] = 8'b10111110;
DRAM[19366] = 8'b11000001;
DRAM[19367] = 8'b11010101;
DRAM[19368] = 8'b11010110;
DRAM[19369] = 8'b11010111;
DRAM[19370] = 8'b11100100;
DRAM[19371] = 8'b11100000;
DRAM[19372] = 8'b11001011;
DRAM[19373] = 8'b11010000;
DRAM[19374] = 8'b11100001;
DRAM[19375] = 8'b11100001;
DRAM[19376] = 8'b11101001;
DRAM[19377] = 8'b11101011;
DRAM[19378] = 8'b11101111;
DRAM[19379] = 8'b11110010;
DRAM[19380] = 8'b11110000;
DRAM[19381] = 8'b11101100;
DRAM[19382] = 8'b11100110;
DRAM[19383] = 8'b11100010;
DRAM[19384] = 8'b11100011;
DRAM[19385] = 8'b11001010;
DRAM[19386] = 8'b11011100;
DRAM[19387] = 8'b11011100;
DRAM[19388] = 8'b10110010;
DRAM[19389] = 8'b10101111;
DRAM[19390] = 8'b10100110;
DRAM[19391] = 8'b1101010;
DRAM[19392] = 8'b1100000;
DRAM[19393] = 8'b1100101;
DRAM[19394] = 8'b10010101;
DRAM[19395] = 8'b10010011;
DRAM[19396] = 8'b10100100;
DRAM[19397] = 8'b11010110;
DRAM[19398] = 8'b11011000;
DRAM[19399] = 8'b11101100;
DRAM[19400] = 8'b11111010;
DRAM[19401] = 8'b11111001;
DRAM[19402] = 8'b11110101;
DRAM[19403] = 8'b11110011;
DRAM[19404] = 8'b11110111;
DRAM[19405] = 8'b11111100;
DRAM[19406] = 8'b11111101;
DRAM[19407] = 8'b11111010;
DRAM[19408] = 8'b11111010;
DRAM[19409] = 8'b11110111;
DRAM[19410] = 8'b11110111;
DRAM[19411] = 8'b11110111;
DRAM[19412] = 8'b11110001;
DRAM[19413] = 8'b11101000;
DRAM[19414] = 8'b11100101;
DRAM[19415] = 8'b11101001;
DRAM[19416] = 8'b11011111;
DRAM[19417] = 8'b11101001;
DRAM[19418] = 8'b11110110;
DRAM[19419] = 8'b11111110;
DRAM[19420] = 8'b11111011;
DRAM[19421] = 8'b11110111;
DRAM[19422] = 8'b11111001;
DRAM[19423] = 8'b11111111;
DRAM[19424] = 8'b11111100;
DRAM[19425] = 8'b11111101;
DRAM[19426] = 8'b11111101;
DRAM[19427] = 8'b11111110;
DRAM[19428] = 8'b11111110;
DRAM[19429] = 8'b11111110;
DRAM[19430] = 8'b11111101;
DRAM[19431] = 8'b11111101;
DRAM[19432] = 8'b11111111;
DRAM[19433] = 8'b11101111;
DRAM[19434] = 8'b10111110;
DRAM[19435] = 8'b10001010;
DRAM[19436] = 8'b1110001;
DRAM[19437] = 8'b1101111;
DRAM[19438] = 8'b1101011;
DRAM[19439] = 8'b1100001;
DRAM[19440] = 8'b1100100;
DRAM[19441] = 8'b1100010;
DRAM[19442] = 8'b1011111;
DRAM[19443] = 8'b1011101;
DRAM[19444] = 8'b1011110;
DRAM[19445] = 8'b1011110;
DRAM[19446] = 8'b1011101;
DRAM[19447] = 8'b1011100;
DRAM[19448] = 8'b1011101;
DRAM[19449] = 8'b1011100;
DRAM[19450] = 8'b1011100;
DRAM[19451] = 8'b1011100;
DRAM[19452] = 8'b1011011;
DRAM[19453] = 8'b1011011;
DRAM[19454] = 8'b1011011;
DRAM[19455] = 8'b1011011;
DRAM[19456] = 8'b1101111;
DRAM[19457] = 8'b1101111;
DRAM[19458] = 8'b1110000;
DRAM[19459] = 8'b1110001;
DRAM[19460] = 8'b1110001;
DRAM[19461] = 8'b1110001;
DRAM[19462] = 8'b1110001;
DRAM[19463] = 8'b1110001;
DRAM[19464] = 8'b1110001;
DRAM[19465] = 8'b1110010;
DRAM[19466] = 8'b1110010;
DRAM[19467] = 8'b1110010;
DRAM[19468] = 8'b1110011;
DRAM[19469] = 8'b1110011;
DRAM[19470] = 8'b1110011;
DRAM[19471] = 8'b1110011;
DRAM[19472] = 8'b1110101;
DRAM[19473] = 8'b1110110;
DRAM[19474] = 8'b1110110;
DRAM[19475] = 8'b1110111;
DRAM[19476] = 8'b1111000;
DRAM[19477] = 8'b1111001;
DRAM[19478] = 8'b1111010;
DRAM[19479] = 8'b1111011;
DRAM[19480] = 8'b1110101;
DRAM[19481] = 8'b1110101;
DRAM[19482] = 8'b1111001;
DRAM[19483] = 8'b1111101;
DRAM[19484] = 8'b10000010;
DRAM[19485] = 8'b10011000;
DRAM[19486] = 8'b11000101;
DRAM[19487] = 8'b11101110;
DRAM[19488] = 8'b11111100;
DRAM[19489] = 8'b11111110;
DRAM[19490] = 8'b11111110;
DRAM[19491] = 8'b11111100;
DRAM[19492] = 8'b11111000;
DRAM[19493] = 8'b11111000;
DRAM[19494] = 8'b11111101;
DRAM[19495] = 8'b11111111;
DRAM[19496] = 8'b11111110;
DRAM[19497] = 8'b11111110;
DRAM[19498] = 8'b11111111;
DRAM[19499] = 8'b11111111;
DRAM[19500] = 8'b11111111;
DRAM[19501] = 8'b11111110;
DRAM[19502] = 8'b11111101;
DRAM[19503] = 8'b11111100;
DRAM[19504] = 8'b11110010;
DRAM[19505] = 8'b11101010;
DRAM[19506] = 8'b11101100;
DRAM[19507] = 8'b11111010;
DRAM[19508] = 8'b11111111;
DRAM[19509] = 8'b11110101;
DRAM[19510] = 8'b11101001;
DRAM[19511] = 8'b11100101;
DRAM[19512] = 8'b11101110;
DRAM[19513] = 8'b11110100;
DRAM[19514] = 8'b11111000;
DRAM[19515] = 8'b11111001;
DRAM[19516] = 8'b11111010;
DRAM[19517] = 8'b11110110;
DRAM[19518] = 8'b11101000;
DRAM[19519] = 8'b11011001;
DRAM[19520] = 8'b11000111;
DRAM[19521] = 8'b11010011;
DRAM[19522] = 8'b11110100;
DRAM[19523] = 8'b11100100;
DRAM[19524] = 8'b11100010;
DRAM[19525] = 8'b11011011;
DRAM[19526] = 8'b11100100;
DRAM[19527] = 8'b11100110;
DRAM[19528] = 8'b11110010;
DRAM[19529] = 8'b10111001;
DRAM[19530] = 8'b11010011;
DRAM[19531] = 8'b10111111;
DRAM[19532] = 8'b10010110;
DRAM[19533] = 8'b10010100;
DRAM[19534] = 8'b1111111;
DRAM[19535] = 8'b1100001;
DRAM[19536] = 8'b1011110;
DRAM[19537] = 8'b1111111;
DRAM[19538] = 8'b10011101;
DRAM[19539] = 8'b10100110;
DRAM[19540] = 8'b10100100;
DRAM[19541] = 8'b10100101;
DRAM[19542] = 8'b10110101;
DRAM[19543] = 8'b11001001;
DRAM[19544] = 8'b11010001;
DRAM[19545] = 8'b11010101;
DRAM[19546] = 8'b11010100;
DRAM[19547] = 8'b11010010;
DRAM[19548] = 8'b11011001;
DRAM[19549] = 8'b11100101;
DRAM[19550] = 8'b11100100;
DRAM[19551] = 8'b11011011;
DRAM[19552] = 8'b11100100;
DRAM[19553] = 8'b11101001;
DRAM[19554] = 8'b11101111;
DRAM[19555] = 8'b11101101;
DRAM[19556] = 8'b11100111;
DRAM[19557] = 8'b11100011;
DRAM[19558] = 8'b11100100;
DRAM[19559] = 8'b11100111;
DRAM[19560] = 8'b11011010;
DRAM[19561] = 8'b11010001;
DRAM[19562] = 8'b11001110;
DRAM[19563] = 8'b11010111;
DRAM[19564] = 8'b11100010;
DRAM[19565] = 8'b11100101;
DRAM[19566] = 8'b11100010;
DRAM[19567] = 8'b11011111;
DRAM[19568] = 8'b11010001;
DRAM[19569] = 8'b11001100;
DRAM[19570] = 8'b11010100;
DRAM[19571] = 8'b11000111;
DRAM[19572] = 8'b10110001;
DRAM[19573] = 8'b11000100;
DRAM[19574] = 8'b10111000;
DRAM[19575] = 8'b11001001;
DRAM[19576] = 8'b11000110;
DRAM[19577] = 8'b10111100;
DRAM[19578] = 8'b11010001;
DRAM[19579] = 8'b10110100;
DRAM[19580] = 8'b10110111;
DRAM[19581] = 8'b11001111;
DRAM[19582] = 8'b10110010;
DRAM[19583] = 8'b10111111;
DRAM[19584] = 8'b11001100;
DRAM[19585] = 8'b11000101;
DRAM[19586] = 8'b11001100;
DRAM[19587] = 8'b11010101;
DRAM[19588] = 8'b11010100;
DRAM[19589] = 8'b11010110;
DRAM[19590] = 8'b11011010;
DRAM[19591] = 8'b11010110;
DRAM[19592] = 8'b11010111;
DRAM[19593] = 8'b11011000;
DRAM[19594] = 8'b11011011;
DRAM[19595] = 8'b11010100;
DRAM[19596] = 8'b11001101;
DRAM[19597] = 8'b11001101;
DRAM[19598] = 8'b11001100;
DRAM[19599] = 8'b11010001;
DRAM[19600] = 8'b11011010;
DRAM[19601] = 8'b11010110;
DRAM[19602] = 8'b11001000;
DRAM[19603] = 8'b10111000;
DRAM[19604] = 8'b10110110;
DRAM[19605] = 8'b11000001;
DRAM[19606] = 8'b11001000;
DRAM[19607] = 8'b11001000;
DRAM[19608] = 8'b10111001;
DRAM[19609] = 8'b10110111;
DRAM[19610] = 8'b10111110;
DRAM[19611] = 8'b10111001;
DRAM[19612] = 8'b10111111;
DRAM[19613] = 8'b11000110;
DRAM[19614] = 8'b10110101;
DRAM[19615] = 8'b10110011;
DRAM[19616] = 8'b11000101;
DRAM[19617] = 8'b11000110;
DRAM[19618] = 8'b10111011;
DRAM[19619] = 8'b10110110;
DRAM[19620] = 8'b10111111;
DRAM[19621] = 8'b11001110;
DRAM[19622] = 8'b11010100;
DRAM[19623] = 8'b11001001;
DRAM[19624] = 8'b11000100;
DRAM[19625] = 8'b11010101;
DRAM[19626] = 8'b11010000;
DRAM[19627] = 8'b11000101;
DRAM[19628] = 8'b11001101;
DRAM[19629] = 8'b11010011;
DRAM[19630] = 8'b11011001;
DRAM[19631] = 8'b11101001;
DRAM[19632] = 8'b11011110;
DRAM[19633] = 8'b11100010;
DRAM[19634] = 8'b11101000;
DRAM[19635] = 8'b11101100;
DRAM[19636] = 8'b11101101;
DRAM[19637] = 8'b11101011;
DRAM[19638] = 8'b11100111;
DRAM[19639] = 8'b11100100;
DRAM[19640] = 8'b11100000;
DRAM[19641] = 8'b11101000;
DRAM[19642] = 8'b11010011;
DRAM[19643] = 8'b10110110;
DRAM[19644] = 8'b10101101;
DRAM[19645] = 8'b10011000;
DRAM[19646] = 8'b1101111;
DRAM[19647] = 8'b1010100;
DRAM[19648] = 8'b110111;
DRAM[19649] = 8'b1001000;
DRAM[19650] = 8'b10010011;
DRAM[19651] = 8'b10011001;
DRAM[19652] = 8'b10010100;
DRAM[19653] = 8'b10110101;
DRAM[19654] = 8'b11000011;
DRAM[19655] = 8'b11100111;
DRAM[19656] = 8'b11110011;
DRAM[19657] = 8'b11111001;
DRAM[19658] = 8'b11111011;
DRAM[19659] = 8'b11110101;
DRAM[19660] = 8'b11110011;
DRAM[19661] = 8'b11110111;
DRAM[19662] = 8'b11111010;
DRAM[19663] = 8'b11111010;
DRAM[19664] = 8'b11111111;
DRAM[19665] = 8'b11111101;
DRAM[19666] = 8'b11111100;
DRAM[19667] = 8'b11111011;
DRAM[19668] = 8'b11110110;
DRAM[19669] = 8'b11110000;
DRAM[19670] = 8'b11101101;
DRAM[19671] = 8'b11101110;
DRAM[19672] = 8'b11100110;
DRAM[19673] = 8'b11100110;
DRAM[19674] = 8'b11101101;
DRAM[19675] = 8'b11110111;
DRAM[19676] = 8'b11111010;
DRAM[19677] = 8'b11111001;
DRAM[19678] = 8'b11111010;
DRAM[19679] = 8'b11111111;
DRAM[19680] = 8'b11111111;
DRAM[19681] = 8'b11111110;
DRAM[19682] = 8'b11111101;
DRAM[19683] = 8'b11111101;
DRAM[19684] = 8'b11111100;
DRAM[19685] = 8'b11111100;
DRAM[19686] = 8'b11111100;
DRAM[19687] = 8'b11111100;
DRAM[19688] = 8'b11111101;
DRAM[19689] = 8'b11111111;
DRAM[19690] = 8'b11101011;
DRAM[19691] = 8'b10111100;
DRAM[19692] = 8'b10010100;
DRAM[19693] = 8'b10000001;
DRAM[19694] = 8'b1110110;
DRAM[19695] = 8'b1101011;
DRAM[19696] = 8'b1101011;
DRAM[19697] = 8'b1100111;
DRAM[19698] = 8'b1100011;
DRAM[19699] = 8'b1100000;
DRAM[19700] = 8'b1011111;
DRAM[19701] = 8'b1011110;
DRAM[19702] = 8'b1011101;
DRAM[19703] = 8'b1011100;
DRAM[19704] = 8'b1011101;
DRAM[19705] = 8'b1011101;
DRAM[19706] = 8'b1011101;
DRAM[19707] = 8'b1011101;
DRAM[19708] = 8'b1011100;
DRAM[19709] = 8'b1011100;
DRAM[19710] = 8'b1011100;
DRAM[19711] = 8'b1011011;
DRAM[19712] = 8'b1101111;
DRAM[19713] = 8'b1110000;
DRAM[19714] = 8'b1110001;
DRAM[19715] = 8'b1110010;
DRAM[19716] = 8'b1110010;
DRAM[19717] = 8'b1110010;
DRAM[19718] = 8'b1110010;
DRAM[19719] = 8'b1110001;
DRAM[19720] = 8'b1110010;
DRAM[19721] = 8'b1110010;
DRAM[19722] = 8'b1110011;
DRAM[19723] = 8'b1110011;
DRAM[19724] = 8'b1110011;
DRAM[19725] = 8'b1110100;
DRAM[19726] = 8'b1110100;
DRAM[19727] = 8'b1110100;
DRAM[19728] = 8'b1110011;
DRAM[19729] = 8'b1110011;
DRAM[19730] = 8'b1110101;
DRAM[19731] = 8'b1110111;
DRAM[19732] = 8'b1111001;
DRAM[19733] = 8'b1111100;
DRAM[19734] = 8'b1111111;
DRAM[19735] = 8'b10000001;
DRAM[19736] = 8'b10000000;
DRAM[19737] = 8'b1111000;
DRAM[19738] = 8'b1110101;
DRAM[19739] = 8'b10000000;
DRAM[19740] = 8'b10011110;
DRAM[19741] = 8'b11000111;
DRAM[19742] = 8'b11101101;
DRAM[19743] = 8'b11111111;
DRAM[19744] = 8'b11111000;
DRAM[19745] = 8'b11111000;
DRAM[19746] = 8'b11111010;
DRAM[19747] = 8'b11111110;
DRAM[19748] = 8'b11111111;
DRAM[19749] = 8'b11111111;
DRAM[19750] = 8'b11111111;
DRAM[19751] = 8'b11111101;
DRAM[19752] = 8'b11111111;
DRAM[19753] = 8'b11111111;
DRAM[19754] = 8'b11111110;
DRAM[19755] = 8'b11111100;
DRAM[19756] = 8'b11111010;
DRAM[19757] = 8'b11110111;
DRAM[19758] = 8'b11110101;
DRAM[19759] = 8'b11110100;
DRAM[19760] = 8'b11101101;
DRAM[19761] = 8'b11110011;
DRAM[19762] = 8'b11111010;
DRAM[19763] = 8'b11111010;
DRAM[19764] = 8'b11101111;
DRAM[19765] = 8'b11100110;
DRAM[19766] = 8'b11100111;
DRAM[19767] = 8'b11101110;
DRAM[19768] = 8'b11110100;
DRAM[19769] = 8'b11111000;
DRAM[19770] = 8'b11111000;
DRAM[19771] = 8'b11110101;
DRAM[19772] = 8'b11110101;
DRAM[19773] = 8'b11110100;
DRAM[19774] = 8'b11101000;
DRAM[19775] = 8'b11011000;
DRAM[19776] = 8'b11010101;
DRAM[19777] = 8'b11011101;
DRAM[19778] = 8'b11110010;
DRAM[19779] = 8'b11011110;
DRAM[19780] = 8'b11011000;
DRAM[19781] = 8'b11010110;
DRAM[19782] = 8'b11101011;
DRAM[19783] = 8'b11100100;
DRAM[19784] = 8'b11100000;
DRAM[19785] = 8'b11000110;
DRAM[19786] = 8'b11000011;
DRAM[19787] = 8'b11000100;
DRAM[19788] = 8'b10100011;
DRAM[19789] = 8'b10001010;
DRAM[19790] = 8'b10000110;
DRAM[19791] = 8'b1010011;
DRAM[19792] = 8'b1001101;
DRAM[19793] = 8'b1100100;
DRAM[19794] = 8'b1111000;
DRAM[19795] = 8'b10010011;
DRAM[19796] = 8'b10110110;
DRAM[19797] = 8'b11000111;
DRAM[19798] = 8'b11000111;
DRAM[19799] = 8'b11001001;
DRAM[19800] = 8'b11010000;
DRAM[19801] = 8'b11010101;
DRAM[19802] = 8'b11011000;
DRAM[19803] = 8'b11011001;
DRAM[19804] = 8'b11011101;
DRAM[19805] = 8'b11100010;
DRAM[19806] = 8'b11100010;
DRAM[19807] = 8'b11011111;
DRAM[19808] = 8'b11011111;
DRAM[19809] = 8'b11100110;
DRAM[19810] = 8'b11101101;
DRAM[19811] = 8'b11101110;
DRAM[19812] = 8'b11101001;
DRAM[19813] = 8'b11100100;
DRAM[19814] = 8'b11100010;
DRAM[19815] = 8'b11100011;
DRAM[19816] = 8'b11011101;
DRAM[19817] = 8'b11010011;
DRAM[19818] = 8'b11001100;
DRAM[19819] = 8'b11001110;
DRAM[19820] = 8'b11010011;
DRAM[19821] = 8'b11010110;
DRAM[19822] = 8'b11011001;
DRAM[19823] = 8'b11011100;
DRAM[19824] = 8'b11010000;
DRAM[19825] = 8'b11001010;
DRAM[19826] = 8'b11001010;
DRAM[19827] = 8'b11010011;
DRAM[19828] = 8'b10110110;
DRAM[19829] = 8'b11000100;
DRAM[19830] = 8'b10111001;
DRAM[19831] = 8'b11000011;
DRAM[19832] = 8'b11000111;
DRAM[19833] = 8'b10111010;
DRAM[19834] = 8'b11001111;
DRAM[19835] = 8'b10111000;
DRAM[19836] = 8'b10110101;
DRAM[19837] = 8'b11001100;
DRAM[19838] = 8'b10111010;
DRAM[19839] = 8'b11000111;
DRAM[19840] = 8'b11000000;
DRAM[19841] = 8'b10111101;
DRAM[19842] = 8'b11001000;
DRAM[19843] = 8'b11010010;
DRAM[19844] = 8'b11001110;
DRAM[19845] = 8'b11001110;
DRAM[19846] = 8'b11010100;
DRAM[19847] = 8'b11010011;
DRAM[19848] = 8'b11010110;
DRAM[19849] = 8'b11010101;
DRAM[19850] = 8'b11011101;
DRAM[19851] = 8'b11010010;
DRAM[19852] = 8'b11001101;
DRAM[19853] = 8'b11010011;
DRAM[19854] = 8'b11001100;
DRAM[19855] = 8'b11010010;
DRAM[19856] = 8'b11011010;
DRAM[19857] = 8'b11010110;
DRAM[19858] = 8'b11000111;
DRAM[19859] = 8'b10110111;
DRAM[19860] = 8'b10110100;
DRAM[19861] = 8'b10111011;
DRAM[19862] = 8'b10111100;
DRAM[19863] = 8'b10110110;
DRAM[19864] = 8'b10101011;
DRAM[19865] = 8'b10110110;
DRAM[19866] = 8'b11000010;
DRAM[19867] = 8'b10111000;
DRAM[19868] = 8'b10111001;
DRAM[19869] = 8'b10111010;
DRAM[19870] = 8'b10101010;
DRAM[19871] = 8'b10110011;
DRAM[19872] = 8'b11000100;
DRAM[19873] = 8'b10111110;
DRAM[19874] = 8'b10101111;
DRAM[19875] = 8'b10111011;
DRAM[19876] = 8'b11000110;
DRAM[19877] = 8'b11000110;
DRAM[19878] = 8'b11001101;
DRAM[19879] = 8'b11000101;
DRAM[19880] = 8'b11001001;
DRAM[19881] = 8'b11010001;
DRAM[19882] = 8'b10111011;
DRAM[19883] = 8'b10110100;
DRAM[19884] = 8'b11010010;
DRAM[19885] = 8'b11011000;
DRAM[19886] = 8'b11001110;
DRAM[19887] = 8'b11011010;
DRAM[19888] = 8'b11011011;
DRAM[19889] = 8'b11011111;
DRAM[19890] = 8'b11100011;
DRAM[19891] = 8'b11100111;
DRAM[19892] = 8'b11101000;
DRAM[19893] = 8'b11100111;
DRAM[19894] = 8'b11100100;
DRAM[19895] = 8'b11100001;
DRAM[19896] = 8'b11100011;
DRAM[19897] = 8'b11010011;
DRAM[19898] = 8'b11011101;
DRAM[19899] = 8'b11011000;
DRAM[19900] = 8'b10110111;
DRAM[19901] = 8'b10101111;
DRAM[19902] = 8'b10011110;
DRAM[19903] = 8'b1101001;
DRAM[19904] = 8'b1001000;
DRAM[19905] = 8'b111010;
DRAM[19906] = 8'b1110111;
DRAM[19907] = 8'b10100010;
DRAM[19908] = 8'b10100100;
DRAM[19909] = 8'b10101100;
DRAM[19910] = 8'b10111100;
DRAM[19911] = 8'b11100010;
DRAM[19912] = 8'b11101101;
DRAM[19913] = 8'b11111001;
DRAM[19914] = 8'b11111111;
DRAM[19915] = 8'b11111000;
DRAM[19916] = 8'b11110011;
DRAM[19917] = 8'b11110101;
DRAM[19918] = 8'b11110111;
DRAM[19919] = 8'b11110101;
DRAM[19920] = 8'b11111001;
DRAM[19921] = 8'b11111010;
DRAM[19922] = 8'b11111011;
DRAM[19923] = 8'b11111010;
DRAM[19924] = 8'b11110101;
DRAM[19925] = 8'b11101100;
DRAM[19926] = 8'b11100010;
DRAM[19927] = 8'b11011101;
DRAM[19928] = 8'b11110011;
DRAM[19929] = 8'b11100001;
DRAM[19930] = 8'b11011000;
DRAM[19931] = 8'b11100101;
DRAM[19932] = 8'b11110111;
DRAM[19933] = 8'b11111110;
DRAM[19934] = 8'b11111101;
DRAM[19935] = 8'b11111100;
DRAM[19936] = 8'b11111111;
DRAM[19937] = 8'b11111111;
DRAM[19938] = 8'b11111101;
DRAM[19939] = 8'b11111011;
DRAM[19940] = 8'b11111010;
DRAM[19941] = 8'b11111010;
DRAM[19942] = 8'b11111010;
DRAM[19943] = 8'b11111011;
DRAM[19944] = 8'b11111001;
DRAM[19945] = 8'b11111111;
DRAM[19946] = 8'b11101111;
DRAM[19947] = 8'b11000000;
DRAM[19948] = 8'b10010001;
DRAM[19949] = 8'b1111010;
DRAM[19950] = 8'b1110100;
DRAM[19951] = 8'b1110010;
DRAM[19952] = 8'b1101101;
DRAM[19953] = 8'b1101001;
DRAM[19954] = 8'b1100100;
DRAM[19955] = 8'b1100001;
DRAM[19956] = 8'b1100000;
DRAM[19957] = 8'b1011111;
DRAM[19958] = 8'b1011111;
DRAM[19959] = 8'b1011110;
DRAM[19960] = 8'b1011110;
DRAM[19961] = 8'b1011110;
DRAM[19962] = 8'b1011110;
DRAM[19963] = 8'b1011101;
DRAM[19964] = 8'b1011101;
DRAM[19965] = 8'b1011101;
DRAM[19966] = 8'b1011100;
DRAM[19967] = 8'b1011100;
DRAM[19968] = 8'b1110000;
DRAM[19969] = 8'b1110001;
DRAM[19970] = 8'b1110001;
DRAM[19971] = 8'b1110010;
DRAM[19972] = 8'b1110011;
DRAM[19973] = 8'b1110011;
DRAM[19974] = 8'b1110010;
DRAM[19975] = 8'b1110010;
DRAM[19976] = 8'b1110011;
DRAM[19977] = 8'b1110011;
DRAM[19978] = 8'b1110011;
DRAM[19979] = 8'b1110100;
DRAM[19980] = 8'b1110100;
DRAM[19981] = 8'b1110100;
DRAM[19982] = 8'b1110101;
DRAM[19983] = 8'b1110101;
DRAM[19984] = 8'b1110100;
DRAM[19985] = 8'b1110100;
DRAM[19986] = 8'b1110101;
DRAM[19987] = 8'b1110111;
DRAM[19988] = 8'b1111010;
DRAM[19989] = 8'b1111101;
DRAM[19990] = 8'b10000000;
DRAM[19991] = 8'b10000010;
DRAM[19992] = 8'b10001011;
DRAM[19993] = 8'b10001010;
DRAM[19994] = 8'b10001100;
DRAM[19995] = 8'b10011011;
DRAM[19996] = 8'b11000000;
DRAM[19997] = 8'b11101000;
DRAM[19998] = 8'b11111001;
DRAM[19999] = 8'b11110111;
DRAM[20000] = 8'b11110110;
DRAM[20001] = 8'b11111000;
DRAM[20002] = 8'b11111011;
DRAM[20003] = 8'b11111111;
DRAM[20004] = 8'b11111111;
DRAM[20005] = 8'b11111111;
DRAM[20006] = 8'b11111101;
DRAM[20007] = 8'b11111010;
DRAM[20008] = 8'b11111110;
DRAM[20009] = 8'b11111110;
DRAM[20010] = 8'b11111101;
DRAM[20011] = 8'b11111011;
DRAM[20012] = 8'b11111000;
DRAM[20013] = 8'b11110101;
DRAM[20014] = 8'b11110011;
DRAM[20015] = 8'b11110001;
DRAM[20016] = 8'b11110101;
DRAM[20017] = 8'b11111000;
DRAM[20018] = 8'b11110010;
DRAM[20019] = 8'b11100101;
DRAM[20020] = 8'b11011100;
DRAM[20021] = 8'b11100001;
DRAM[20022] = 8'b11110000;
DRAM[20023] = 8'b11111011;
DRAM[20024] = 8'b11110110;
DRAM[20025] = 8'b11111000;
DRAM[20026] = 8'b11110101;
DRAM[20027] = 8'b11101111;
DRAM[20028] = 8'b11110000;
DRAM[20029] = 8'b11110010;
DRAM[20030] = 8'b11101000;
DRAM[20031] = 8'b11011000;
DRAM[20032] = 8'b11100101;
DRAM[20033] = 8'b11100101;
DRAM[20034] = 8'b11101111;
DRAM[20035] = 8'b11011110;
DRAM[20036] = 8'b11011011;
DRAM[20037] = 8'b11011111;
DRAM[20038] = 8'b11110110;
DRAM[20039] = 8'b11100001;
DRAM[20040] = 8'b11010101;
DRAM[20041] = 8'b11001011;
DRAM[20042] = 8'b10110000;
DRAM[20043] = 8'b11001001;
DRAM[20044] = 8'b10011011;
DRAM[20045] = 8'b10011011;
DRAM[20046] = 8'b1110001;
DRAM[20047] = 8'b1001011;
DRAM[20048] = 8'b111111;
DRAM[20049] = 8'b1101001;
DRAM[20050] = 8'b10000110;
DRAM[20051] = 8'b10010010;
DRAM[20052] = 8'b10100010;
DRAM[20053] = 8'b10101011;
DRAM[20054] = 8'b10110111;
DRAM[20055] = 8'b11001110;
DRAM[20056] = 8'b11001110;
DRAM[20057] = 8'b11010101;
DRAM[20058] = 8'b11011101;
DRAM[20059] = 8'b11100001;
DRAM[20060] = 8'b11011101;
DRAM[20061] = 8'b11011010;
DRAM[20062] = 8'b11100001;
DRAM[20063] = 8'b11101011;
DRAM[20064] = 8'b11100010;
DRAM[20065] = 8'b11100111;
DRAM[20066] = 8'b11101100;
DRAM[20067] = 8'b11101101;
DRAM[20068] = 8'b11101001;
DRAM[20069] = 8'b11100100;
DRAM[20070] = 8'b11100001;
DRAM[20071] = 8'b11100000;
DRAM[20072] = 8'b11101010;
DRAM[20073] = 8'b11011111;
DRAM[20074] = 8'b11010011;
DRAM[20075] = 8'b11001011;
DRAM[20076] = 8'b11000110;
DRAM[20077] = 8'b11000110;
DRAM[20078] = 8'b11001110;
DRAM[20079] = 8'b11011000;
DRAM[20080] = 8'b11010011;
DRAM[20081] = 8'b11000101;
DRAM[20082] = 8'b11000010;
DRAM[20083] = 8'b11010101;
DRAM[20084] = 8'b11000101;
DRAM[20085] = 8'b10111011;
DRAM[20086] = 8'b11000100;
DRAM[20087] = 8'b10111111;
DRAM[20088] = 8'b11000111;
DRAM[20089] = 8'b10110111;
DRAM[20090] = 8'b11000011;
DRAM[20091] = 8'b10110111;
DRAM[20092] = 8'b10110011;
DRAM[20093] = 8'b11000100;
DRAM[20094] = 8'b10111110;
DRAM[20095] = 8'b11000110;
DRAM[20096] = 8'b10110101;
DRAM[20097] = 8'b10110110;
DRAM[20098] = 8'b11000101;
DRAM[20099] = 8'b11001101;
DRAM[20100] = 8'b11000100;
DRAM[20101] = 8'b11000011;
DRAM[20102] = 8'b11001110;
DRAM[20103] = 8'b11010011;
DRAM[20104] = 8'b11010010;
DRAM[20105] = 8'b11001111;
DRAM[20106] = 8'b11011100;
DRAM[20107] = 8'b11001111;
DRAM[20108] = 8'b11001100;
DRAM[20109] = 8'b11011000;
DRAM[20110] = 8'b11001110;
DRAM[20111] = 8'b11010101;
DRAM[20112] = 8'b11010110;
DRAM[20113] = 8'b11010011;
DRAM[20114] = 8'b11000111;
DRAM[20115] = 8'b10111010;
DRAM[20116] = 8'b10110111;
DRAM[20117] = 8'b10111011;
DRAM[20118] = 8'b10110110;
DRAM[20119] = 8'b10101100;
DRAM[20120] = 8'b10011110;
DRAM[20121] = 8'b10110110;
DRAM[20122] = 8'b11000101;
DRAM[20123] = 8'b10110011;
DRAM[20124] = 8'b10101100;
DRAM[20125] = 8'b10101010;
DRAM[20126] = 8'b10100110;
DRAM[20127] = 8'b11000001;
DRAM[20128] = 8'b11000010;
DRAM[20129] = 8'b10110011;
DRAM[20130] = 8'b10101000;
DRAM[20131] = 8'b11001011;
DRAM[20132] = 8'b11010010;
DRAM[20133] = 8'b10111001;
DRAM[20134] = 8'b11000011;
DRAM[20135] = 8'b11001101;
DRAM[20136] = 8'b11010010;
DRAM[20137] = 8'b11001011;
DRAM[20138] = 8'b11000001;
DRAM[20139] = 8'b11000011;
DRAM[20140] = 8'b11001111;
DRAM[20141] = 8'b11010010;
DRAM[20142] = 8'b11001110;
DRAM[20143] = 8'b11001110;
DRAM[20144] = 8'b11011110;
DRAM[20145] = 8'b11100000;
DRAM[20146] = 8'b11100010;
DRAM[20147] = 8'b11100100;
DRAM[20148] = 8'b11100011;
DRAM[20149] = 8'b11100001;
DRAM[20150] = 8'b11011110;
DRAM[20151] = 8'b11011100;
DRAM[20152] = 8'b11100111;
DRAM[20153] = 8'b11110111;
DRAM[20154] = 8'b11100110;
DRAM[20155] = 8'b11010100;
DRAM[20156] = 8'b11010011;
DRAM[20157] = 8'b10110100;
DRAM[20158] = 8'b10000110;
DRAM[20159] = 8'b1111001;
DRAM[20160] = 8'b1110001;
DRAM[20161] = 8'b1000011;
DRAM[20162] = 8'b1011000;
DRAM[20163] = 8'b10010100;
DRAM[20164] = 8'b10101011;
DRAM[20165] = 8'b10110101;
DRAM[20166] = 8'b11000110;
DRAM[20167] = 8'b11010000;
DRAM[20168] = 8'b11101100;
DRAM[20169] = 8'b11111001;
DRAM[20170] = 8'b11111111;
DRAM[20171] = 8'b11111010;
DRAM[20172] = 8'b11110110;
DRAM[20173] = 8'b11110111;
DRAM[20174] = 8'b11110100;
DRAM[20175] = 8'b11101101;
DRAM[20176] = 8'b11101100;
DRAM[20177] = 8'b11101111;
DRAM[20178] = 8'b11110001;
DRAM[20179] = 8'b11110001;
DRAM[20180] = 8'b11101110;
DRAM[20181] = 8'b11100111;
DRAM[20182] = 8'b11011101;
DRAM[20183] = 8'b11010110;
DRAM[20184] = 8'b11100110;
DRAM[20185] = 8'b11010111;
DRAM[20186] = 8'b11010010;
DRAM[20187] = 8'b11100010;
DRAM[20188] = 8'b11110011;
DRAM[20189] = 8'b11111001;
DRAM[20190] = 8'b11111001;
DRAM[20191] = 8'b11111100;
DRAM[20192] = 8'b11111111;
DRAM[20193] = 8'b11111101;
DRAM[20194] = 8'b11111011;
DRAM[20195] = 8'b11111000;
DRAM[20196] = 8'b11111000;
DRAM[20197] = 8'b11111000;
DRAM[20198] = 8'b11111010;
DRAM[20199] = 8'b11111011;
DRAM[20200] = 8'b11111101;
DRAM[20201] = 8'b11111001;
DRAM[20202] = 8'b11100001;
DRAM[20203] = 8'b10110110;
DRAM[20204] = 8'b10001101;
DRAM[20205] = 8'b1110110;
DRAM[20206] = 8'b1110000;
DRAM[20207] = 8'b1101111;
DRAM[20208] = 8'b1101011;
DRAM[20209] = 8'b1100111;
DRAM[20210] = 8'b1100011;
DRAM[20211] = 8'b1100000;
DRAM[20212] = 8'b1100000;
DRAM[20213] = 8'b1100001;
DRAM[20214] = 8'b1100001;
DRAM[20215] = 8'b1100001;
DRAM[20216] = 8'b1011111;
DRAM[20217] = 8'b1011111;
DRAM[20218] = 8'b1011110;
DRAM[20219] = 8'b1011110;
DRAM[20220] = 8'b1011110;
DRAM[20221] = 8'b1011101;
DRAM[20222] = 8'b1011101;
DRAM[20223] = 8'b1011101;
DRAM[20224] = 8'b1110000;
DRAM[20225] = 8'b1110001;
DRAM[20226] = 8'b1110010;
DRAM[20227] = 8'b1110011;
DRAM[20228] = 8'b1110011;
DRAM[20229] = 8'b1110011;
DRAM[20230] = 8'b1110011;
DRAM[20231] = 8'b1110010;
DRAM[20232] = 8'b1110011;
DRAM[20233] = 8'b1110011;
DRAM[20234] = 8'b1110100;
DRAM[20235] = 8'b1110100;
DRAM[20236] = 8'b1110100;
DRAM[20237] = 8'b1110101;
DRAM[20238] = 8'b1110101;
DRAM[20239] = 8'b1110101;
DRAM[20240] = 8'b1111000;
DRAM[20241] = 8'b1111000;
DRAM[20242] = 8'b1110111;
DRAM[20243] = 8'b1111000;
DRAM[20244] = 8'b1111001;
DRAM[20245] = 8'b1111100;
DRAM[20246] = 8'b1111110;
DRAM[20247] = 8'b1111111;
DRAM[20248] = 8'b10001001;
DRAM[20249] = 8'b10011011;
DRAM[20250] = 8'b10101100;
DRAM[20251] = 8'b10111100;
DRAM[20252] = 8'b11011010;
DRAM[20253] = 8'b11111010;
DRAM[20254] = 8'b11111111;
DRAM[20255] = 8'b11110110;
DRAM[20256] = 8'b11111111;
DRAM[20257] = 8'b11111111;
DRAM[20258] = 8'b11111110;
DRAM[20259] = 8'b11111011;
DRAM[20260] = 8'b11111000;
DRAM[20261] = 8'b11111000;
DRAM[20262] = 8'b11111010;
DRAM[20263] = 8'b11111100;
DRAM[20264] = 8'b11111100;
DRAM[20265] = 8'b11111100;
DRAM[20266] = 8'b11111100;
DRAM[20267] = 8'b11111011;
DRAM[20268] = 8'b11111010;
DRAM[20269] = 8'b11111001;
DRAM[20270] = 8'b11110111;
DRAM[20271] = 8'b11110110;
DRAM[20272] = 8'b11111000;
DRAM[20273] = 8'b11110100;
DRAM[20274] = 8'b11101000;
DRAM[20275] = 8'b11100000;
DRAM[20276] = 8'b11100111;
DRAM[20277] = 8'b11110111;
DRAM[20278] = 8'b11111100;
DRAM[20279] = 8'b11110110;
DRAM[20280] = 8'b11110110;
DRAM[20281] = 8'b11111000;
DRAM[20282] = 8'b11110011;
DRAM[20283] = 8'b11101001;
DRAM[20284] = 8'b11100110;
DRAM[20285] = 8'b11100101;
DRAM[20286] = 8'b11010111;
DRAM[20287] = 8'b11000100;
DRAM[20288] = 8'b11100011;
DRAM[20289] = 8'b11100000;
DRAM[20290] = 8'b11101000;
DRAM[20291] = 8'b11011101;
DRAM[20292] = 8'b11100010;
DRAM[20293] = 8'b11100111;
DRAM[20294] = 8'b11111001;
DRAM[20295] = 8'b11010110;
DRAM[20296] = 8'b11011101;
DRAM[20297] = 8'b10110010;
DRAM[20298] = 8'b11000110;
DRAM[20299] = 8'b10101011;
DRAM[20300] = 8'b10100011;
DRAM[20301] = 8'b10100010;
DRAM[20302] = 8'b1011100;
DRAM[20303] = 8'b1000100;
DRAM[20304] = 8'b1010111;
DRAM[20305] = 8'b1110101;
DRAM[20306] = 8'b10000001;
DRAM[20307] = 8'b10000111;
DRAM[20308] = 8'b10011101;
DRAM[20309] = 8'b10100101;
DRAM[20310] = 8'b10101000;
DRAM[20311] = 8'b10110111;
DRAM[20312] = 8'b11001100;
DRAM[20313] = 8'b11000001;
DRAM[20314] = 8'b11000001;
DRAM[20315] = 8'b11010010;
DRAM[20316] = 8'b11100011;
DRAM[20317] = 8'b11100111;
DRAM[20318] = 8'b11101000;
DRAM[20319] = 8'b11101010;
DRAM[20320] = 8'b11011011;
DRAM[20321] = 8'b11011111;
DRAM[20322] = 8'b11100100;
DRAM[20323] = 8'b11100110;
DRAM[20324] = 8'b11100110;
DRAM[20325] = 8'b11100101;
DRAM[20326] = 8'b11100011;
DRAM[20327] = 8'b11100011;
DRAM[20328] = 8'b11011100;
DRAM[20329] = 8'b11011100;
DRAM[20330] = 8'b11011101;
DRAM[20331] = 8'b11011011;
DRAM[20332] = 8'b11010010;
DRAM[20333] = 8'b11001010;
DRAM[20334] = 8'b11001010;
DRAM[20335] = 8'b11010000;
DRAM[20336] = 8'b11011001;
DRAM[20337] = 8'b11000010;
DRAM[20338] = 8'b11000000;
DRAM[20339] = 8'b11010001;
DRAM[20340] = 8'b11010010;
DRAM[20341] = 8'b10110001;
DRAM[20342] = 8'b11001101;
DRAM[20343] = 8'b10111100;
DRAM[20344] = 8'b11001100;
DRAM[20345] = 8'b10111000;
DRAM[20346] = 8'b10111011;
DRAM[20347] = 8'b10111000;
DRAM[20348] = 8'b10110101;
DRAM[20349] = 8'b11000000;
DRAM[20350] = 8'b11000001;
DRAM[20351] = 8'b11000100;
DRAM[20352] = 8'b10101111;
DRAM[20353] = 8'b10110010;
DRAM[20354] = 8'b11000010;
DRAM[20355] = 8'b11001000;
DRAM[20356] = 8'b10111100;
DRAM[20357] = 8'b10111100;
DRAM[20358] = 8'b11001011;
DRAM[20359] = 8'b11010100;
DRAM[20360] = 8'b11001011;
DRAM[20361] = 8'b11001001;
DRAM[20362] = 8'b11011001;
DRAM[20363] = 8'b11001011;
DRAM[20364] = 8'b11001010;
DRAM[20365] = 8'b11011001;
DRAM[20366] = 8'b11001110;
DRAM[20367] = 8'b11010101;
DRAM[20368] = 8'b11010000;
DRAM[20369] = 8'b11001111;
DRAM[20370] = 8'b11000111;
DRAM[20371] = 8'b10111101;
DRAM[20372] = 8'b10111101;
DRAM[20373] = 8'b11000001;
DRAM[20374] = 8'b10111001;
DRAM[20375] = 8'b10101101;
DRAM[20376] = 8'b10110010;
DRAM[20377] = 8'b10111010;
DRAM[20378] = 8'b10111000;
DRAM[20379] = 8'b10100101;
DRAM[20380] = 8'b10101110;
DRAM[20381] = 8'b10110111;
DRAM[20382] = 8'b10110010;
DRAM[20383] = 8'b11001010;
DRAM[20384] = 8'b10110011;
DRAM[20385] = 8'b11000011;
DRAM[20386] = 8'b10111101;
DRAM[20387] = 8'b11001101;
DRAM[20388] = 8'b11010001;
DRAM[20389] = 8'b11001001;
DRAM[20390] = 8'b11010111;
DRAM[20391] = 8'b11001101;
DRAM[20392] = 8'b11001010;
DRAM[20393] = 8'b10111110;
DRAM[20394] = 8'b11010000;
DRAM[20395] = 8'b11011100;
DRAM[20396] = 8'b11001010;
DRAM[20397] = 8'b11001011;
DRAM[20398] = 8'b11011100;
DRAM[20399] = 8'b11011001;
DRAM[20400] = 8'b11011001;
DRAM[20401] = 8'b11011010;
DRAM[20402] = 8'b11011101;
DRAM[20403] = 8'b11100000;
DRAM[20404] = 8'b11100010;
DRAM[20405] = 8'b11100010;
DRAM[20406] = 8'b11100001;
DRAM[20407] = 8'b11100000;
DRAM[20408] = 8'b11011101;
DRAM[20409] = 8'b11011101;
DRAM[20410] = 8'b11001101;
DRAM[20411] = 8'b11000001;
DRAM[20412] = 8'b11000001;
DRAM[20413] = 8'b10110110;
DRAM[20414] = 8'b10100110;
DRAM[20415] = 8'b10100010;
DRAM[20416] = 8'b1110010;
DRAM[20417] = 8'b1001110;
DRAM[20418] = 8'b1001111;
DRAM[20419] = 8'b1111100;
DRAM[20420] = 8'b10010000;
DRAM[20421] = 8'b10100111;
DRAM[20422] = 8'b11000111;
DRAM[20423] = 8'b10111111;
DRAM[20424] = 8'b11101101;
DRAM[20425] = 8'b11111000;
DRAM[20426] = 8'b11111101;
DRAM[20427] = 8'b11111010;
DRAM[20428] = 8'b11111001;
DRAM[20429] = 8'b11111011;
DRAM[20430] = 8'b11110011;
DRAM[20431] = 8'b11100101;
DRAM[20432] = 8'b11100111;
DRAM[20433] = 8'b11101000;
DRAM[20434] = 8'b11101010;
DRAM[20435] = 8'b11101010;
DRAM[20436] = 8'b11101011;
DRAM[20437] = 8'b11101011;
DRAM[20438] = 8'b11101000;
DRAM[20439] = 8'b11100100;
DRAM[20440] = 8'b11001010;
DRAM[20441] = 8'b11001110;
DRAM[20442] = 8'b11011100;
DRAM[20443] = 8'b11101100;
DRAM[20444] = 8'b11110000;
DRAM[20445] = 8'b11101100;
DRAM[20446] = 8'b11110001;
DRAM[20447] = 8'b11111101;
DRAM[20448] = 8'b11111101;
DRAM[20449] = 8'b11111011;
DRAM[20450] = 8'b11111001;
DRAM[20451] = 8'b11110111;
DRAM[20452] = 8'b11110111;
DRAM[20453] = 8'b11111000;
DRAM[20454] = 8'b11111011;
DRAM[20455] = 8'b11111101;
DRAM[20456] = 8'b11111111;
DRAM[20457] = 8'b11111010;
DRAM[20458] = 8'b11101011;
DRAM[20459] = 8'b11010000;
DRAM[20460] = 8'b10110000;
DRAM[20461] = 8'b10010001;
DRAM[20462] = 8'b1111000;
DRAM[20463] = 8'b1101010;
DRAM[20464] = 8'b1101000;
DRAM[20465] = 8'b1100100;
DRAM[20466] = 8'b1100000;
DRAM[20467] = 8'b1011110;
DRAM[20468] = 8'b1011111;
DRAM[20469] = 8'b1100010;
DRAM[20470] = 8'b1100011;
DRAM[20471] = 8'b1100011;
DRAM[20472] = 8'b1011111;
DRAM[20473] = 8'b1011111;
DRAM[20474] = 8'b1011111;
DRAM[20475] = 8'b1011110;
DRAM[20476] = 8'b1011110;
DRAM[20477] = 8'b1011110;
DRAM[20478] = 8'b1011101;
DRAM[20479] = 8'b1011101;
DRAM[20480] = 8'b1110010;
DRAM[20481] = 8'b1110010;
DRAM[20482] = 8'b1110010;
DRAM[20483] = 8'b1110011;
DRAM[20484] = 8'b1110011;
DRAM[20485] = 8'b1110100;
DRAM[20486] = 8'b1110100;
DRAM[20487] = 8'b1110100;
DRAM[20488] = 8'b1110110;
DRAM[20489] = 8'b1110110;
DRAM[20490] = 8'b1110110;
DRAM[20491] = 8'b1110111;
DRAM[20492] = 8'b1110111;
DRAM[20493] = 8'b1110111;
DRAM[20494] = 8'b1111000;
DRAM[20495] = 8'b1111000;
DRAM[20496] = 8'b1110101;
DRAM[20497] = 8'b1111000;
DRAM[20498] = 8'b1111100;
DRAM[20499] = 8'b1111101;
DRAM[20500] = 8'b1111100;
DRAM[20501] = 8'b1111010;
DRAM[20502] = 8'b1111001;
DRAM[20503] = 8'b1111001;
DRAM[20504] = 8'b10000101;
DRAM[20505] = 8'b10000100;
DRAM[20506] = 8'b10001100;
DRAM[20507] = 8'b10101001;
DRAM[20508] = 8'b11011001;
DRAM[20509] = 8'b11111111;
DRAM[20510] = 8'b11111111;
DRAM[20511] = 8'b11111010;
DRAM[20512] = 8'b11111010;
DRAM[20513] = 8'b11111001;
DRAM[20514] = 8'b11111001;
DRAM[20515] = 8'b11111010;
DRAM[20516] = 8'b11111100;
DRAM[20517] = 8'b11111110;
DRAM[20518] = 8'b11111111;
DRAM[20519] = 8'b11111111;
DRAM[20520] = 8'b11111001;
DRAM[20521] = 8'b11111110;
DRAM[20522] = 8'b11111101;
DRAM[20523] = 8'b11110101;
DRAM[20524] = 8'b11110011;
DRAM[20525] = 8'b11111001;
DRAM[20526] = 8'b11111101;
DRAM[20527] = 8'b11111011;
DRAM[20528] = 8'b11110000;
DRAM[20529] = 8'b11100111;
DRAM[20530] = 8'b11101101;
DRAM[20531] = 8'b11010101;
DRAM[20532] = 8'b11011011;
DRAM[20533] = 8'b11111001;
DRAM[20534] = 8'b11110000;
DRAM[20535] = 8'b11110100;
DRAM[20536] = 8'b11111111;
DRAM[20537] = 8'b11110100;
DRAM[20538] = 8'b11010000;
DRAM[20539] = 8'b11011000;
DRAM[20540] = 8'b11111011;
DRAM[20541] = 8'b11011100;
DRAM[20542] = 8'b10111010;
DRAM[20543] = 8'b11011000;
DRAM[20544] = 8'b11100100;
DRAM[20545] = 8'b11110100;
DRAM[20546] = 8'b11101101;
DRAM[20547] = 8'b11001011;
DRAM[20548] = 8'b11101011;
DRAM[20549] = 8'b11001110;
DRAM[20550] = 8'b11101111;
DRAM[20551] = 8'b11100111;
DRAM[20552] = 8'b11000111;
DRAM[20553] = 8'b11001001;
DRAM[20554] = 8'b10111110;
DRAM[20555] = 8'b10111010;
DRAM[20556] = 8'b10011000;
DRAM[20557] = 8'b10001101;
DRAM[20558] = 8'b1100001;
DRAM[20559] = 8'b111100;
DRAM[20560] = 8'b1100101;
DRAM[20561] = 8'b1110011;
DRAM[20562] = 8'b10000011;
DRAM[20563] = 8'b10001111;
DRAM[20564] = 8'b10010110;
DRAM[20565] = 8'b10100001;
DRAM[20566] = 8'b10110010;
DRAM[20567] = 8'b10111111;
DRAM[20568] = 8'b11000010;
DRAM[20569] = 8'b11010011;
DRAM[20570] = 8'b11100010;
DRAM[20571] = 8'b11011110;
DRAM[20572] = 8'b11001101;
DRAM[20573] = 8'b11000010;
DRAM[20574] = 8'b11001000;
DRAM[20575] = 8'b11010011;
DRAM[20576] = 8'b11101110;
DRAM[20577] = 8'b11100100;
DRAM[20578] = 8'b11011010;
DRAM[20579] = 8'b11011000;
DRAM[20580] = 8'b11011011;
DRAM[20581] = 8'b11011011;
DRAM[20582] = 8'b11010101;
DRAM[20583] = 8'b11001101;
DRAM[20584] = 8'b11000100;
DRAM[20585] = 8'b11001100;
DRAM[20586] = 8'b11010101;
DRAM[20587] = 8'b11011001;
DRAM[20588] = 8'b11010100;
DRAM[20589] = 8'b11001101;
DRAM[20590] = 8'b11001000;
DRAM[20591] = 8'b11000110;
DRAM[20592] = 8'b11010001;
DRAM[20593] = 8'b11010110;
DRAM[20594] = 8'b11010010;
DRAM[20595] = 8'b11000111;
DRAM[20596] = 8'b11000111;
DRAM[20597] = 8'b11001101;
DRAM[20598] = 8'b11000101;
DRAM[20599] = 8'b10110100;
DRAM[20600] = 8'b11001001;
DRAM[20601] = 8'b11000011;
DRAM[20602] = 8'b10101010;
DRAM[20603] = 8'b11000000;
DRAM[20604] = 8'b11000111;
DRAM[20605] = 8'b10101101;
DRAM[20606] = 8'b10111010;
DRAM[20607] = 8'b11000110;
DRAM[20608] = 8'b10110110;
DRAM[20609] = 8'b10101011;
DRAM[20610] = 8'b11000111;
DRAM[20611] = 8'b11001001;
DRAM[20612] = 8'b11000011;
DRAM[20613] = 8'b11001001;
DRAM[20614] = 8'b11000001;
DRAM[20615] = 8'b11001100;
DRAM[20616] = 8'b11001100;
DRAM[20617] = 8'b11001010;
DRAM[20618] = 8'b11001100;
DRAM[20619] = 8'b11001011;
DRAM[20620] = 8'b11001010;
DRAM[20621] = 8'b11010011;
DRAM[20622] = 8'b11010100;
DRAM[20623] = 8'b11000101;
DRAM[20624] = 8'b11010001;
DRAM[20625] = 8'b11001001;
DRAM[20626] = 8'b10111100;
DRAM[20627] = 8'b10111010;
DRAM[20628] = 8'b11000010;
DRAM[20629] = 8'b10111000;
DRAM[20630] = 8'b10100111;
DRAM[20631] = 8'b10100011;
DRAM[20632] = 8'b10101110;
DRAM[20633] = 8'b10110001;
DRAM[20634] = 8'b10110111;
DRAM[20635] = 8'b10110101;
DRAM[20636] = 8'b10110001;
DRAM[20637] = 8'b10111010;
DRAM[20638] = 8'b10111111;
DRAM[20639] = 8'b10110101;
DRAM[20640] = 8'b10101010;
DRAM[20641] = 8'b10111100;
DRAM[20642] = 8'b11000110;
DRAM[20643] = 8'b11001011;
DRAM[20644] = 8'b11010100;
DRAM[20645] = 8'b11010000;
DRAM[20646] = 8'b11000011;
DRAM[20647] = 8'b10111111;
DRAM[20648] = 8'b10111110;
DRAM[20649] = 8'b11001000;
DRAM[20650] = 8'b11010100;
DRAM[20651] = 8'b11011010;
DRAM[20652] = 8'b11010111;
DRAM[20653] = 8'b11010010;
DRAM[20654] = 8'b11010000;
DRAM[20655] = 8'b11010000;
DRAM[20656] = 8'b11010001;
DRAM[20657] = 8'b11010110;
DRAM[20658] = 8'b11011111;
DRAM[20659] = 8'b11101001;
DRAM[20660] = 8'b11110000;
DRAM[20661] = 8'b11110001;
DRAM[20662] = 8'b11101101;
DRAM[20663] = 8'b11101001;
DRAM[20664] = 8'b11100011;
DRAM[20665] = 8'b11011110;
DRAM[20666] = 8'b11011001;
DRAM[20667] = 8'b11011010;
DRAM[20668] = 8'b11010111;
DRAM[20669] = 8'b11000111;
DRAM[20670] = 8'b10101010;
DRAM[20671] = 8'b10010000;
DRAM[20672] = 8'b10001101;
DRAM[20673] = 8'b1110111;
DRAM[20674] = 8'b10000110;
DRAM[20675] = 8'b10000010;
DRAM[20676] = 8'b10011011;
DRAM[20677] = 8'b10111011;
DRAM[20678] = 8'b11011111;
DRAM[20679] = 8'b11000010;
DRAM[20680] = 8'b11110001;
DRAM[20681] = 8'b11111010;
DRAM[20682] = 8'b11111100;
DRAM[20683] = 8'b11111001;
DRAM[20684] = 8'b11111011;
DRAM[20685] = 8'b11111101;
DRAM[20686] = 8'b11110010;
DRAM[20687] = 8'b11100011;
DRAM[20688] = 8'b11001011;
DRAM[20689] = 8'b11110111;
DRAM[20690] = 8'b11011100;
DRAM[20691] = 8'b11110101;
DRAM[20692] = 8'b11011101;
DRAM[20693] = 8'b11110001;
DRAM[20694] = 8'b11100110;
DRAM[20695] = 8'b11100000;
DRAM[20696] = 8'b11011010;
DRAM[20697] = 8'b10110010;
DRAM[20698] = 8'b11011101;
DRAM[20699] = 8'b11011000;
DRAM[20700] = 8'b11011101;
DRAM[20701] = 8'b11110000;
DRAM[20702] = 8'b11111111;
DRAM[20703] = 8'b11101101;
DRAM[20704] = 8'b11111110;
DRAM[20705] = 8'b11110010;
DRAM[20706] = 8'b11111001;
DRAM[20707] = 8'b11111000;
DRAM[20708] = 8'b11101001;
DRAM[20709] = 8'b11110101;
DRAM[20710] = 8'b11111111;
DRAM[20711] = 8'b11110000;
DRAM[20712] = 8'b11111111;
DRAM[20713] = 8'b11110001;
DRAM[20714] = 8'b11110011;
DRAM[20715] = 8'b10101101;
DRAM[20716] = 8'b10011000;
DRAM[20717] = 8'b10010110;
DRAM[20718] = 8'b10000101;
DRAM[20719] = 8'b1101010;
DRAM[20720] = 8'b1100110;
DRAM[20721] = 8'b1100100;
DRAM[20722] = 8'b1100011;
DRAM[20723] = 8'b1100011;
DRAM[20724] = 8'b1100011;
DRAM[20725] = 8'b1100011;
DRAM[20726] = 8'b1100001;
DRAM[20727] = 8'b1100000;
DRAM[20728] = 8'b1011111;
DRAM[20729] = 8'b1011111;
DRAM[20730] = 8'b1011111;
DRAM[20731] = 8'b1011111;
DRAM[20732] = 8'b1011111;
DRAM[20733] = 8'b1011111;
DRAM[20734] = 8'b1011111;
DRAM[20735] = 8'b1011111;
DRAM[20736] = 8'b1110010;
DRAM[20737] = 8'b1110010;
DRAM[20738] = 8'b1110010;
DRAM[20739] = 8'b1110011;
DRAM[20740] = 8'b1110011;
DRAM[20741] = 8'b1110011;
DRAM[20742] = 8'b1110100;
DRAM[20743] = 8'b1110100;
DRAM[20744] = 8'b1110110;
DRAM[20745] = 8'b1110110;
DRAM[20746] = 8'b1110111;
DRAM[20747] = 8'b1110111;
DRAM[20748] = 8'b1110111;
DRAM[20749] = 8'b1111000;
DRAM[20750] = 8'b1111000;
DRAM[20751] = 8'b1111000;
DRAM[20752] = 8'b1111001;
DRAM[20753] = 8'b1111010;
DRAM[20754] = 8'b1111010;
DRAM[20755] = 8'b1111010;
DRAM[20756] = 8'b1111010;
DRAM[20757] = 8'b1111011;
DRAM[20758] = 8'b1111110;
DRAM[20759] = 8'b10000001;
DRAM[20760] = 8'b10000011;
DRAM[20761] = 8'b1101010;
DRAM[20762] = 8'b1111110;
DRAM[20763] = 8'b11000110;
DRAM[20764] = 8'b11111010;
DRAM[20765] = 8'b11111100;
DRAM[20766] = 8'b11110101;
DRAM[20767] = 8'b11111101;
DRAM[20768] = 8'b11111011;
DRAM[20769] = 8'b11111010;
DRAM[20770] = 8'b11111011;
DRAM[20771] = 8'b11111100;
DRAM[20772] = 8'b11111110;
DRAM[20773] = 8'b11111110;
DRAM[20774] = 8'b11111110;
DRAM[20775] = 8'b11111101;
DRAM[20776] = 8'b11111001;
DRAM[20777] = 8'b11111010;
DRAM[20778] = 8'b11111010;
DRAM[20779] = 8'b11111001;
DRAM[20780] = 8'b11111010;
DRAM[20781] = 8'b11111000;
DRAM[20782] = 8'b11110010;
DRAM[20783] = 8'b11101011;
DRAM[20784] = 8'b11110000;
DRAM[20785] = 8'b11011101;
DRAM[20786] = 8'b11001110;
DRAM[20787] = 8'b11011110;
DRAM[20788] = 8'b11110000;
DRAM[20789] = 8'b11110010;
DRAM[20790] = 8'b11101111;
DRAM[20791] = 8'b11100111;
DRAM[20792] = 8'b11110010;
DRAM[20793] = 8'b11100110;
DRAM[20794] = 8'b11100100;
DRAM[20795] = 8'b11110011;
DRAM[20796] = 8'b11101111;
DRAM[20797] = 8'b11001111;
DRAM[20798] = 8'b11001100;
DRAM[20799] = 8'b11101110;
DRAM[20800] = 8'b11011001;
DRAM[20801] = 8'b11110010;
DRAM[20802] = 8'b11010110;
DRAM[20803] = 8'b11100100;
DRAM[20804] = 8'b11011100;
DRAM[20805] = 8'b11101100;
DRAM[20806] = 8'b11101001;
DRAM[20807] = 8'b11100010;
DRAM[20808] = 8'b11001000;
DRAM[20809] = 8'b11001010;
DRAM[20810] = 8'b10110010;
DRAM[20811] = 8'b10110110;
DRAM[20812] = 8'b10010111;
DRAM[20813] = 8'b10001101;
DRAM[20814] = 8'b1011101;
DRAM[20815] = 8'b1000111;
DRAM[20816] = 8'b1100100;
DRAM[20817] = 8'b1101101;
DRAM[20818] = 8'b1111100;
DRAM[20819] = 8'b10001100;
DRAM[20820] = 8'b10100000;
DRAM[20821] = 8'b10110111;
DRAM[20822] = 8'b11001111;
DRAM[20823] = 8'b11011111;
DRAM[20824] = 8'b11011010;
DRAM[20825] = 8'b11010101;
DRAM[20826] = 8'b11001111;
DRAM[20827] = 8'b11001111;
DRAM[20828] = 8'b11010010;
DRAM[20829] = 8'b11010100;
DRAM[20830] = 8'b11010001;
DRAM[20831] = 8'b11001110;
DRAM[20832] = 8'b11001101;
DRAM[20833] = 8'b11010011;
DRAM[20834] = 8'b11011010;
DRAM[20835] = 8'b11011111;
DRAM[20836] = 8'b11011110;
DRAM[20837] = 8'b11010111;
DRAM[20838] = 8'b11001100;
DRAM[20839] = 8'b11000101;
DRAM[20840] = 8'b11001000;
DRAM[20841] = 8'b11000111;
DRAM[20842] = 8'b11001000;
DRAM[20843] = 8'b11001110;
DRAM[20844] = 8'b11010011;
DRAM[20845] = 8'b11010000;
DRAM[20846] = 8'b11000101;
DRAM[20847] = 8'b10111011;
DRAM[20848] = 8'b11000101;
DRAM[20849] = 8'b11001010;
DRAM[20850] = 8'b11001001;
DRAM[20851] = 8'b11000100;
DRAM[20852] = 8'b11000101;
DRAM[20853] = 8'b11001101;
DRAM[20854] = 8'b11001110;
DRAM[20855] = 8'b11001000;
DRAM[20856] = 8'b10110101;
DRAM[20857] = 8'b11000000;
DRAM[20858] = 8'b10111010;
DRAM[20859] = 8'b10111100;
DRAM[20860] = 8'b10111001;
DRAM[20861] = 8'b10101010;
DRAM[20862] = 8'b10110101;
DRAM[20863] = 8'b11000110;
DRAM[20864] = 8'b10110011;
DRAM[20865] = 8'b10101100;
DRAM[20866] = 8'b11000111;
DRAM[20867] = 8'b11001011;
DRAM[20868] = 8'b11000010;
DRAM[20869] = 8'b11000101;
DRAM[20870] = 8'b10111101;
DRAM[20871] = 8'b11000101;
DRAM[20872] = 8'b11000001;
DRAM[20873] = 8'b11001001;
DRAM[20874] = 8'b11001001;
DRAM[20875] = 8'b11000101;
DRAM[20876] = 8'b11000111;
DRAM[20877] = 8'b11001110;
DRAM[20878] = 8'b11001110;
DRAM[20879] = 8'b11001001;
DRAM[20880] = 8'b11001011;
DRAM[20881] = 8'b11001000;
DRAM[20882] = 8'b10111101;
DRAM[20883] = 8'b10111011;
DRAM[20884] = 8'b10111110;
DRAM[20885] = 8'b10110010;
DRAM[20886] = 8'b10100010;
DRAM[20887] = 8'b10100001;
DRAM[20888] = 8'b10110111;
DRAM[20889] = 8'b10111011;
DRAM[20890] = 8'b10110110;
DRAM[20891] = 8'b10101111;
DRAM[20892] = 8'b10110010;
DRAM[20893] = 8'b10111001;
DRAM[20894] = 8'b10111000;
DRAM[20895] = 8'b10110011;
DRAM[20896] = 8'b10111010;
DRAM[20897] = 8'b11001010;
DRAM[20898] = 8'b11001101;
DRAM[20899] = 8'b11001001;
DRAM[20900] = 8'b11001001;
DRAM[20901] = 8'b11000011;
DRAM[20902] = 8'b10111011;
DRAM[20903] = 8'b10111100;
DRAM[20904] = 8'b11010000;
DRAM[20905] = 8'b11010010;
DRAM[20906] = 8'b11010100;
DRAM[20907] = 8'b11010010;
DRAM[20908] = 8'b11001100;
DRAM[20909] = 8'b11000100;
DRAM[20910] = 8'b10111100;
DRAM[20911] = 8'b10110111;
DRAM[20912] = 8'b11010000;
DRAM[20913] = 8'b11010011;
DRAM[20914] = 8'b11010111;
DRAM[20915] = 8'b11011100;
DRAM[20916] = 8'b11011111;
DRAM[20917] = 8'b11011111;
DRAM[20918] = 8'b11011101;
DRAM[20919] = 8'b11011011;
DRAM[20920] = 8'b11011001;
DRAM[20921] = 8'b11011001;
DRAM[20922] = 8'b11010101;
DRAM[20923] = 8'b11010001;
DRAM[20924] = 8'b11001110;
DRAM[20925] = 8'b11001000;
DRAM[20926] = 8'b10110110;
DRAM[20927] = 8'b10100100;
DRAM[20928] = 8'b10010001;
DRAM[20929] = 8'b1101010;
DRAM[20930] = 8'b1111010;
DRAM[20931] = 8'b10000110;
DRAM[20932] = 8'b10101000;
DRAM[20933] = 8'b10011111;
DRAM[20934] = 8'b10111001;
DRAM[20935] = 8'b10110110;
DRAM[20936] = 8'b11011101;
DRAM[20937] = 8'b11110010;
DRAM[20938] = 8'b11111001;
DRAM[20939] = 8'b11110100;
DRAM[20940] = 8'b11110101;
DRAM[20941] = 8'b11110100;
DRAM[20942] = 8'b11101101;
DRAM[20943] = 8'b11101011;
DRAM[20944] = 8'b11001111;
DRAM[20945] = 8'b11011100;
DRAM[20946] = 8'b11011110;
DRAM[20947] = 8'b11011101;
DRAM[20948] = 8'b11100110;
DRAM[20949] = 8'b11011100;
DRAM[20950] = 8'b11101111;
DRAM[20951] = 8'b11011110;
DRAM[20952] = 8'b11011000;
DRAM[20953] = 8'b11100101;
DRAM[20954] = 8'b11001110;
DRAM[20955] = 8'b11011110;
DRAM[20956] = 8'b11100001;
DRAM[20957] = 8'b11101001;
DRAM[20958] = 8'b11100000;
DRAM[20959] = 8'b11110010;
DRAM[20960] = 8'b11110110;
DRAM[20961] = 8'b11110111;
DRAM[20962] = 8'b11111000;
DRAM[20963] = 8'b11111011;
DRAM[20964] = 8'b11110111;
DRAM[20965] = 8'b11101001;
DRAM[20966] = 8'b11101010;
DRAM[20967] = 8'b11111010;
DRAM[20968] = 8'b11111100;
DRAM[20969] = 8'b11110011;
DRAM[20970] = 8'b11100011;
DRAM[20971] = 8'b10100111;
DRAM[20972] = 8'b10000111;
DRAM[20973] = 8'b10000001;
DRAM[20974] = 8'b1111010;
DRAM[20975] = 8'b1101000;
DRAM[20976] = 8'b1100111;
DRAM[20977] = 8'b1100101;
DRAM[20978] = 8'b1100011;
DRAM[20979] = 8'b1100011;
DRAM[20980] = 8'b1100100;
DRAM[20981] = 8'b1100011;
DRAM[20982] = 8'b1100010;
DRAM[20983] = 8'b1100000;
DRAM[20984] = 8'b1011111;
DRAM[20985] = 8'b1011111;
DRAM[20986] = 8'b1011111;
DRAM[20987] = 8'b1011111;
DRAM[20988] = 8'b1011111;
DRAM[20989] = 8'b1011111;
DRAM[20990] = 8'b1011111;
DRAM[20991] = 8'b1011111;
DRAM[20992] = 8'b1110010;
DRAM[20993] = 8'b1110010;
DRAM[20994] = 8'b1110010;
DRAM[20995] = 8'b1110011;
DRAM[20996] = 8'b1110011;
DRAM[20997] = 8'b1110011;
DRAM[20998] = 8'b1110100;
DRAM[20999] = 8'b1110100;
DRAM[21000] = 8'b1110111;
DRAM[21001] = 8'b1110111;
DRAM[21002] = 8'b1110111;
DRAM[21003] = 8'b1111000;
DRAM[21004] = 8'b1111000;
DRAM[21005] = 8'b1111000;
DRAM[21006] = 8'b1111001;
DRAM[21007] = 8'b1111001;
DRAM[21008] = 8'b1111000;
DRAM[21009] = 8'b1111010;
DRAM[21010] = 8'b1111011;
DRAM[21011] = 8'b1111011;
DRAM[21012] = 8'b1111011;
DRAM[21013] = 8'b1111011;
DRAM[21014] = 8'b1111110;
DRAM[21015] = 8'b10000000;
DRAM[21016] = 8'b10000010;
DRAM[21017] = 8'b10001100;
DRAM[21018] = 8'b10110011;
DRAM[21019] = 8'b11101000;
DRAM[21020] = 8'b11111111;
DRAM[21021] = 8'b11111001;
DRAM[21022] = 8'b11110110;
DRAM[21023] = 8'b11111111;
DRAM[21024] = 8'b11111101;
DRAM[21025] = 8'b11111100;
DRAM[21026] = 8'b11111011;
DRAM[21027] = 8'b11111101;
DRAM[21028] = 8'b11111110;
DRAM[21029] = 8'b11111110;
DRAM[21030] = 8'b11111100;
DRAM[21031] = 8'b11111010;
DRAM[21032] = 8'b11111011;
DRAM[21033] = 8'b11110111;
DRAM[21034] = 8'b11110110;
DRAM[21035] = 8'b11111010;
DRAM[21036] = 8'b11111011;
DRAM[21037] = 8'b11110001;
DRAM[21038] = 8'b11100010;
DRAM[21039] = 8'b11011000;
DRAM[21040] = 8'b11010011;
DRAM[21041] = 8'b11011110;
DRAM[21042] = 8'b11010011;
DRAM[21043] = 8'b11101111;
DRAM[21044] = 8'b11110111;
DRAM[21045] = 8'b11101001;
DRAM[21046] = 8'b11111011;
DRAM[21047] = 8'b11110010;
DRAM[21048] = 8'b11100011;
DRAM[21049] = 8'b11100000;
DRAM[21050] = 8'b11110101;
DRAM[21051] = 8'b11111010;
DRAM[21052] = 8'b11011101;
DRAM[21053] = 8'b11010001;
DRAM[21054] = 8'b11100011;
DRAM[21055] = 8'b11101110;
DRAM[21056] = 8'b11011010;
DRAM[21057] = 8'b11101100;
DRAM[21058] = 8'b11010100;
DRAM[21059] = 8'b11110100;
DRAM[21060] = 8'b11011101;
DRAM[21061] = 8'b11111110;
DRAM[21062] = 8'b11101010;
DRAM[21063] = 8'b11010111;
DRAM[21064] = 8'b11010000;
DRAM[21065] = 8'b11010000;
DRAM[21066] = 8'b10101000;
DRAM[21067] = 8'b10110001;
DRAM[21068] = 8'b10010000;
DRAM[21069] = 8'b1111110;
DRAM[21070] = 8'b1000101;
DRAM[21071] = 8'b1001000;
DRAM[21072] = 8'b1011111;
DRAM[21073] = 8'b1101011;
DRAM[21074] = 8'b10000000;
DRAM[21075] = 8'b10010111;
DRAM[21076] = 8'b10101100;
DRAM[21077] = 8'b10111100;
DRAM[21078] = 8'b11000111;
DRAM[21079] = 8'b11001101;
DRAM[21080] = 8'b11010001;
DRAM[21081] = 8'b11010100;
DRAM[21082] = 8'b11011010;
DRAM[21083] = 8'b11011110;
DRAM[21084] = 8'b11011110;
DRAM[21085] = 8'b11011001;
DRAM[21086] = 8'b11010010;
DRAM[21087] = 8'b11001101;
DRAM[21088] = 8'b11001100;
DRAM[21089] = 8'b11000100;
DRAM[21090] = 8'b10111111;
DRAM[21091] = 8'b11000011;
DRAM[21092] = 8'b11001100;
DRAM[21093] = 8'b11001111;
DRAM[21094] = 8'b11001001;
DRAM[21095] = 8'b11000010;
DRAM[21096] = 8'b11000101;
DRAM[21097] = 8'b11000010;
DRAM[21098] = 8'b11000001;
DRAM[21099] = 8'b11000100;
DRAM[21100] = 8'b11001001;
DRAM[21101] = 8'b11001011;
DRAM[21102] = 8'b11000111;
DRAM[21103] = 8'b11000011;
DRAM[21104] = 8'b11000000;
DRAM[21105] = 8'b11000010;
DRAM[21106] = 8'b11000010;
DRAM[21107] = 8'b10111110;
DRAM[21108] = 8'b10111011;
DRAM[21109] = 8'b10111101;
DRAM[21110] = 8'b11000100;
DRAM[21111] = 8'b11001011;
DRAM[21112] = 8'b10111011;
DRAM[21113] = 8'b10111011;
DRAM[21114] = 8'b10111001;
DRAM[21115] = 8'b10101111;
DRAM[21116] = 8'b10111000;
DRAM[21117] = 8'b11000000;
DRAM[21118] = 8'b10110010;
DRAM[21119] = 8'b10110100;
DRAM[21120] = 8'b10110001;
DRAM[21121] = 8'b10101101;
DRAM[21122] = 8'b11000100;
DRAM[21123] = 8'b11001011;
DRAM[21124] = 8'b11000100;
DRAM[21125] = 8'b11000011;
DRAM[21126] = 8'b10111010;
DRAM[21127] = 8'b10111010;
DRAM[21128] = 8'b10111011;
DRAM[21129] = 8'b11001101;
DRAM[21130] = 8'b11001000;
DRAM[21131] = 8'b10111110;
DRAM[21132] = 8'b11000111;
DRAM[21133] = 8'b11001001;
DRAM[21134] = 8'b11000011;
DRAM[21135] = 8'b11001010;
DRAM[21136] = 8'b11000010;
DRAM[21137] = 8'b11000100;
DRAM[21138] = 8'b10111111;
DRAM[21139] = 8'b10111010;
DRAM[21140] = 8'b10111000;
DRAM[21141] = 8'b10101001;
DRAM[21142] = 8'b10011110;
DRAM[21143] = 8'b10100010;
DRAM[21144] = 8'b10111010;
DRAM[21145] = 8'b11000011;
DRAM[21146] = 8'b10110110;
DRAM[21147] = 8'b10101011;
DRAM[21148] = 8'b10111001;
DRAM[21149] = 8'b10111010;
DRAM[21150] = 8'b10101100;
DRAM[21151] = 8'b10101001;
DRAM[21152] = 8'b10110100;
DRAM[21153] = 8'b11000010;
DRAM[21154] = 8'b11000011;
DRAM[21155] = 8'b10111101;
DRAM[21156] = 8'b11000001;
DRAM[21157] = 8'b11000011;
DRAM[21158] = 8'b11000111;
DRAM[21159] = 8'b11010000;
DRAM[21160] = 8'b11100000;
DRAM[21161] = 8'b11010101;
DRAM[21162] = 8'b11000111;
DRAM[21163] = 8'b10111110;
DRAM[21164] = 8'b10111111;
DRAM[21165] = 8'b11000111;
DRAM[21166] = 8'b11001111;
DRAM[21167] = 8'b11010100;
DRAM[21168] = 8'b11001100;
DRAM[21169] = 8'b11001110;
DRAM[21170] = 8'b11010001;
DRAM[21171] = 8'b11010011;
DRAM[21172] = 8'b11010101;
DRAM[21173] = 8'b11010111;
DRAM[21174] = 8'b11011010;
DRAM[21175] = 8'b11011100;
DRAM[21176] = 8'b11100000;
DRAM[21177] = 8'b11100111;
DRAM[21178] = 8'b11100011;
DRAM[21179] = 8'b11010110;
DRAM[21180] = 8'b11001101;
DRAM[21181] = 8'b11000111;
DRAM[21182] = 8'b10110111;
DRAM[21183] = 8'b10100100;
DRAM[21184] = 8'b10010000;
DRAM[21185] = 8'b1011111;
DRAM[21186] = 8'b1010100;
DRAM[21187] = 8'b1011110;
DRAM[21188] = 8'b10001100;
DRAM[21189] = 8'b10000011;
DRAM[21190] = 8'b10100111;
DRAM[21191] = 8'b11001100;
DRAM[21192] = 8'b11001011;
DRAM[21193] = 8'b11101111;
DRAM[21194] = 8'b11111100;
DRAM[21195] = 8'b11110111;
DRAM[21196] = 8'b11111001;
DRAM[21197] = 8'b11110011;
DRAM[21198] = 8'b11101110;
DRAM[21199] = 8'b11111010;
DRAM[21200] = 8'b11001100;
DRAM[21201] = 8'b11000110;
DRAM[21202] = 8'b11011100;
DRAM[21203] = 8'b11011000;
DRAM[21204] = 8'b11011011;
DRAM[21205] = 8'b11000101;
DRAM[21206] = 8'b11101011;
DRAM[21207] = 8'b11100010;
DRAM[21208] = 8'b11011101;
DRAM[21209] = 8'b11011100;
DRAM[21210] = 8'b11000111;
DRAM[21211] = 8'b11101110;
DRAM[21212] = 8'b11011001;
DRAM[21213] = 8'b11011010;
DRAM[21214] = 8'b11110010;
DRAM[21215] = 8'b11101110;
DRAM[21216] = 8'b11101001;
DRAM[21217] = 8'b11111100;
DRAM[21218] = 8'b11110100;
DRAM[21219] = 8'b11110000;
DRAM[21220] = 8'b11111111;
DRAM[21221] = 8'b11110001;
DRAM[21222] = 8'b11100010;
DRAM[21223] = 8'b11110110;
DRAM[21224] = 8'b11111000;
DRAM[21225] = 8'b11110111;
DRAM[21226] = 8'b11001111;
DRAM[21227] = 8'b10100111;
DRAM[21228] = 8'b1111100;
DRAM[21229] = 8'b1110010;
DRAM[21230] = 8'b1110101;
DRAM[21231] = 8'b1101111;
DRAM[21232] = 8'b1100111;
DRAM[21233] = 8'b1100101;
DRAM[21234] = 8'b1100100;
DRAM[21235] = 8'b1100011;
DRAM[21236] = 8'b1100100;
DRAM[21237] = 8'b1100100;
DRAM[21238] = 8'b1100010;
DRAM[21239] = 8'b1100001;
DRAM[21240] = 8'b1100000;
DRAM[21241] = 8'b1100000;
DRAM[21242] = 8'b1100000;
DRAM[21243] = 8'b1100000;
DRAM[21244] = 8'b1100000;
DRAM[21245] = 8'b1100000;
DRAM[21246] = 8'b1100000;
DRAM[21247] = 8'b1100000;
DRAM[21248] = 8'b1110010;
DRAM[21249] = 8'b1110010;
DRAM[21250] = 8'b1110011;
DRAM[21251] = 8'b1110011;
DRAM[21252] = 8'b1110011;
DRAM[21253] = 8'b1110100;
DRAM[21254] = 8'b1110100;
DRAM[21255] = 8'b1110100;
DRAM[21256] = 8'b1111000;
DRAM[21257] = 8'b1111000;
DRAM[21258] = 8'b1111000;
DRAM[21259] = 8'b1111000;
DRAM[21260] = 8'b1111001;
DRAM[21261] = 8'b1111001;
DRAM[21262] = 8'b1111001;
DRAM[21263] = 8'b1111010;
DRAM[21264] = 8'b1110101;
DRAM[21265] = 8'b1111001;
DRAM[21266] = 8'b1111110;
DRAM[21267] = 8'b1111111;
DRAM[21268] = 8'b1111110;
DRAM[21269] = 8'b1111100;
DRAM[21270] = 8'b1111011;
DRAM[21271] = 8'b1111010;
DRAM[21272] = 8'b10010010;
DRAM[21273] = 8'b10110010;
DRAM[21274] = 8'b11011010;
DRAM[21275] = 8'b11110011;
DRAM[21276] = 8'b11111000;
DRAM[21277] = 8'b11110111;
DRAM[21278] = 8'b11111011;
DRAM[21279] = 8'b11111111;
DRAM[21280] = 8'b11111111;
DRAM[21281] = 8'b11111101;
DRAM[21282] = 8'b11111010;
DRAM[21283] = 8'b11111010;
DRAM[21284] = 8'b11111011;
DRAM[21285] = 8'b11111100;
DRAM[21286] = 8'b11111011;
DRAM[21287] = 8'b11111001;
DRAM[21288] = 8'b11111100;
DRAM[21289] = 8'b11110100;
DRAM[21290] = 8'b11110000;
DRAM[21291] = 8'b11110011;
DRAM[21292] = 8'b11110000;
DRAM[21293] = 8'b11100101;
DRAM[21294] = 8'b11011010;
DRAM[21295] = 8'b11010110;
DRAM[21296] = 8'b11000110;
DRAM[21297] = 8'b11101000;
DRAM[21298] = 8'b11101101;
DRAM[21299] = 8'b11101101;
DRAM[21300] = 8'b11101100;
DRAM[21301] = 8'b11110000;
DRAM[21302] = 8'b11111100;
DRAM[21303] = 8'b11101011;
DRAM[21304] = 8'b11011111;
DRAM[21305] = 8'b11101000;
DRAM[21306] = 8'b11110000;
DRAM[21307] = 8'b11100100;
DRAM[21308] = 8'b11010110;
DRAM[21309] = 8'b11100010;
DRAM[21310] = 8'b11101010;
DRAM[21311] = 8'b11011010;
DRAM[21312] = 8'b11100110;
DRAM[21313] = 8'b11100100;
DRAM[21314] = 8'b11101110;
DRAM[21315] = 8'b11101110;
DRAM[21316] = 8'b11110001;
DRAM[21317] = 8'b11110110;
DRAM[21318] = 8'b11110011;
DRAM[21319] = 8'b11001011;
DRAM[21320] = 8'b11010000;
DRAM[21321] = 8'b11010011;
DRAM[21322] = 8'b10100110;
DRAM[21323] = 8'b10110010;
DRAM[21324] = 8'b10001101;
DRAM[21325] = 8'b1110001;
DRAM[21326] = 8'b111000;
DRAM[21327] = 8'b1010001;
DRAM[21328] = 8'b1101101;
DRAM[21329] = 8'b1111100;
DRAM[21330] = 8'b10010001;
DRAM[21331] = 8'b10100011;
DRAM[21332] = 8'b10101111;
DRAM[21333] = 8'b10110101;
DRAM[21334] = 8'b10111000;
DRAM[21335] = 8'b10111001;
DRAM[21336] = 8'b11001001;
DRAM[21337] = 8'b11010011;
DRAM[21338] = 8'b11100000;
DRAM[21339] = 8'b11100110;
DRAM[21340] = 8'b11100010;
DRAM[21341] = 8'b11011011;
DRAM[21342] = 8'b11010110;
DRAM[21343] = 8'b11010100;
DRAM[21344] = 8'b11001101;
DRAM[21345] = 8'b11010010;
DRAM[21346] = 8'b11010010;
DRAM[21347] = 8'b11000111;
DRAM[21348] = 8'b10111010;
DRAM[21349] = 8'b10111011;
DRAM[21350] = 8'b11001011;
DRAM[21351] = 8'b11011100;
DRAM[21352] = 8'b11000100;
DRAM[21353] = 8'b11001010;
DRAM[21354] = 8'b11001100;
DRAM[21355] = 8'b11000110;
DRAM[21356] = 8'b10111101;
DRAM[21357] = 8'b10111010;
DRAM[21358] = 8'b11000000;
DRAM[21359] = 8'b11001000;
DRAM[21360] = 8'b10111100;
DRAM[21361] = 8'b10111101;
DRAM[21362] = 8'b11000000;
DRAM[21363] = 8'b10111110;
DRAM[21364] = 8'b10110110;
DRAM[21365] = 8'b10110001;
DRAM[21366] = 8'b10111001;
DRAM[21367] = 8'b11000110;
DRAM[21368] = 8'b11001000;
DRAM[21369] = 8'b10111001;
DRAM[21370] = 8'b10111000;
DRAM[21371] = 8'b10101011;
DRAM[21372] = 8'b10111100;
DRAM[21373] = 8'b11001011;
DRAM[21374] = 8'b10101111;
DRAM[21375] = 8'b10101111;
DRAM[21376] = 8'b10110001;
DRAM[21377] = 8'b10101100;
DRAM[21378] = 8'b10111011;
DRAM[21379] = 8'b11000110;
DRAM[21380] = 8'b11000111;
DRAM[21381] = 8'b11000111;
DRAM[21382] = 8'b10111101;
DRAM[21383] = 8'b10101111;
DRAM[21384] = 8'b10111111;
DRAM[21385] = 8'b11010011;
DRAM[21386] = 8'b11000110;
DRAM[21387] = 8'b10111000;
DRAM[21388] = 8'b11001000;
DRAM[21389] = 8'b11000111;
DRAM[21390] = 8'b10111010;
DRAM[21391] = 8'b11000011;
DRAM[21392] = 8'b10111010;
DRAM[21393] = 8'b11000000;
DRAM[21394] = 8'b10111100;
DRAM[21395] = 8'b10110110;
DRAM[21396] = 8'b10110001;
DRAM[21397] = 8'b10100100;
DRAM[21398] = 8'b10011111;
DRAM[21399] = 8'b10101010;
DRAM[21400] = 8'b10110011;
DRAM[21401] = 8'b11000011;
DRAM[21402] = 8'b10110100;
DRAM[21403] = 8'b10101010;
DRAM[21404] = 8'b10111110;
DRAM[21405] = 8'b10111010;
DRAM[21406] = 8'b10100010;
DRAM[21407] = 8'b10100001;
DRAM[21408] = 8'b10110110;
DRAM[21409] = 8'b10111110;
DRAM[21410] = 8'b10111010;
DRAM[21411] = 8'b10110100;
DRAM[21412] = 8'b10111110;
DRAM[21413] = 8'b11000110;
DRAM[21414] = 8'b11001100;
DRAM[21415] = 8'b11010110;
DRAM[21416] = 8'b11000010;
DRAM[21417] = 8'b11001000;
DRAM[21418] = 8'b11010000;
DRAM[21419] = 8'b11010111;
DRAM[21420] = 8'b11011010;
DRAM[21421] = 8'b11010111;
DRAM[21422] = 8'b11010001;
DRAM[21423] = 8'b11001100;
DRAM[21424] = 8'b11001000;
DRAM[21425] = 8'b11001011;
DRAM[21426] = 8'b11010001;
DRAM[21427] = 8'b11010101;
DRAM[21428] = 8'b11011001;
DRAM[21429] = 8'b11011110;
DRAM[21430] = 8'b11100100;
DRAM[21431] = 8'b11101001;
DRAM[21432] = 8'b11010111;
DRAM[21433] = 8'b11100001;
DRAM[21434] = 8'b11100000;
DRAM[21435] = 8'b11010001;
DRAM[21436] = 8'b11000101;
DRAM[21437] = 8'b10111100;
DRAM[21438] = 8'b10100100;
DRAM[21439] = 8'b10001010;
DRAM[21440] = 8'b1101100;
DRAM[21441] = 8'b1011011;
DRAM[21442] = 8'b1000110;
DRAM[21443] = 8'b1011110;
DRAM[21444] = 8'b10001000;
DRAM[21445] = 8'b10010001;
DRAM[21446] = 8'b10011100;
DRAM[21447] = 8'b11000101;
DRAM[21448] = 8'b10111110;
DRAM[21449] = 8'b11101000;
DRAM[21450] = 8'b11111011;
DRAM[21451] = 8'b11111100;
DRAM[21452] = 8'b11111111;
DRAM[21453] = 8'b11110110;
DRAM[21454] = 8'b11101110;
DRAM[21455] = 8'b11111101;
DRAM[21456] = 8'b11001110;
DRAM[21457] = 8'b11000001;
DRAM[21458] = 8'b11010101;
DRAM[21459] = 8'b11100110;
DRAM[21460] = 8'b11001000;
DRAM[21461] = 8'b10111110;
DRAM[21462] = 8'b11011001;
DRAM[21463] = 8'b11100101;
DRAM[21464] = 8'b11011101;
DRAM[21465] = 8'b10111110;
DRAM[21466] = 8'b11001100;
DRAM[21467] = 8'b11011111;
DRAM[21468] = 8'b11100000;
DRAM[21469] = 8'b11010000;
DRAM[21470] = 8'b11111000;
DRAM[21471] = 8'b11101000;
DRAM[21472] = 8'b11011111;
DRAM[21473] = 8'b11110111;
DRAM[21474] = 8'b11110000;
DRAM[21475] = 8'b11100000;
DRAM[21476] = 8'b11110010;
DRAM[21477] = 8'b11111111;
DRAM[21478] = 8'b11110110;
DRAM[21479] = 8'b11100110;
DRAM[21480] = 8'b11110100;
DRAM[21481] = 8'b11111000;
DRAM[21482] = 8'b10111101;
DRAM[21483] = 8'b10100111;
DRAM[21484] = 8'b1111100;
DRAM[21485] = 8'b1110000;
DRAM[21486] = 8'b1110100;
DRAM[21487] = 8'b1110101;
DRAM[21488] = 8'b1101000;
DRAM[21489] = 8'b1100110;
DRAM[21490] = 8'b1100100;
DRAM[21491] = 8'b1100100;
DRAM[21492] = 8'b1100101;
DRAM[21493] = 8'b1100101;
DRAM[21494] = 8'b1100011;
DRAM[21495] = 8'b1100001;
DRAM[21496] = 8'b1100001;
DRAM[21497] = 8'b1100001;
DRAM[21498] = 8'b1100001;
DRAM[21499] = 8'b1100001;
DRAM[21500] = 8'b1100000;
DRAM[21501] = 8'b1100000;
DRAM[21502] = 8'b1100000;
DRAM[21503] = 8'b1100000;
DRAM[21504] = 8'b1110011;
DRAM[21505] = 8'b1110100;
DRAM[21506] = 8'b1110100;
DRAM[21507] = 8'b1110100;
DRAM[21508] = 8'b1110101;
DRAM[21509] = 8'b1110101;
DRAM[21510] = 8'b1110101;
DRAM[21511] = 8'b1110110;
DRAM[21512] = 8'b1111000;
DRAM[21513] = 8'b1111001;
DRAM[21514] = 8'b1111001;
DRAM[21515] = 8'b1111001;
DRAM[21516] = 8'b1111010;
DRAM[21517] = 8'b1111010;
DRAM[21518] = 8'b1111010;
DRAM[21519] = 8'b1111010;
DRAM[21520] = 8'b1111000;
DRAM[21521] = 8'b1111010;
DRAM[21522] = 8'b1111100;
DRAM[21523] = 8'b1111110;
DRAM[21524] = 8'b1111110;
DRAM[21525] = 8'b10000000;
DRAM[21526] = 8'b10000011;
DRAM[21527] = 8'b10000101;
DRAM[21528] = 8'b10100110;
DRAM[21529] = 8'b10101011;
DRAM[21530] = 8'b11000110;
DRAM[21531] = 8'b11101101;
DRAM[21532] = 8'b11111111;
DRAM[21533] = 8'b11111010;
DRAM[21534] = 8'b11110111;
DRAM[21535] = 8'b11111111;
DRAM[21536] = 8'b11111111;
DRAM[21537] = 8'b11111101;
DRAM[21538] = 8'b11110110;
DRAM[21539] = 8'b11110100;
DRAM[21540] = 8'b11110110;
DRAM[21541] = 8'b11111001;
DRAM[21542] = 8'b11111001;
DRAM[21543] = 8'b11110111;
DRAM[21544] = 8'b11110100;
DRAM[21545] = 8'b11101110;
DRAM[21546] = 8'b11101001;
DRAM[21547] = 8'b11100101;
DRAM[21548] = 8'b11100001;
DRAM[21549] = 8'b11011110;
DRAM[21550] = 8'b11011111;
DRAM[21551] = 8'b11100100;
DRAM[21552] = 8'b11011111;
DRAM[21553] = 8'b11100100;
DRAM[21554] = 8'b11101111;
DRAM[21555] = 8'b11011111;
DRAM[21556] = 8'b11100110;
DRAM[21557] = 8'b11111011;
DRAM[21558] = 8'b11100101;
DRAM[21559] = 8'b11010011;
DRAM[21560] = 8'b11100001;
DRAM[21561] = 8'b11101001;
DRAM[21562] = 8'b11011111;
DRAM[21563] = 8'b11010110;
DRAM[21564] = 8'b11100000;
DRAM[21565] = 8'b11100100;
DRAM[21566] = 8'b11011101;
DRAM[21567] = 8'b11011100;
DRAM[21568] = 8'b11101001;
DRAM[21569] = 8'b11100001;
DRAM[21570] = 8'b11111110;
DRAM[21571] = 8'b11100110;
DRAM[21572] = 8'b11110101;
DRAM[21573] = 8'b11101101;
DRAM[21574] = 8'b11110011;
DRAM[21575] = 8'b11001001;
DRAM[21576] = 8'b11000110;
DRAM[21577] = 8'b11001001;
DRAM[21578] = 8'b10100111;
DRAM[21579] = 8'b10110011;
DRAM[21580] = 8'b10010001;
DRAM[21581] = 8'b1101100;
DRAM[21582] = 8'b1000000;
DRAM[21583] = 8'b1100111;
DRAM[21584] = 8'b10000100;
DRAM[21585] = 8'b10001110;
DRAM[21586] = 8'b10011100;
DRAM[21587] = 8'b10100101;
DRAM[21588] = 8'b10101011;
DRAM[21589] = 8'b10110101;
DRAM[21590] = 8'b11000100;
DRAM[21591] = 8'b11010000;
DRAM[21592] = 8'b11011001;
DRAM[21593] = 8'b11010010;
DRAM[21594] = 8'b11001100;
DRAM[21595] = 8'b11010000;
DRAM[21596] = 8'b11011001;
DRAM[21597] = 8'b11100000;
DRAM[21598] = 8'b11011111;
DRAM[21599] = 8'b11011010;
DRAM[21600] = 8'b11010010;
DRAM[21601] = 8'b11001101;
DRAM[21602] = 8'b11001000;
DRAM[21603] = 8'b11001000;
DRAM[21604] = 8'b11001011;
DRAM[21605] = 8'b11001000;
DRAM[21606] = 8'b11000000;
DRAM[21607] = 8'b10111000;
DRAM[21608] = 8'b11000100;
DRAM[21609] = 8'b11001010;
DRAM[21610] = 8'b11001111;
DRAM[21611] = 8'b11001011;
DRAM[21612] = 8'b11000000;
DRAM[21613] = 8'b10110111;
DRAM[21614] = 8'b10110101;
DRAM[21615] = 8'b10110111;
DRAM[21616] = 8'b10110101;
DRAM[21617] = 8'b10111000;
DRAM[21618] = 8'b10111110;
DRAM[21619] = 8'b10111111;
DRAM[21620] = 8'b10111000;
DRAM[21621] = 8'b10110010;
DRAM[21622] = 8'b10110111;
DRAM[21623] = 8'b11000010;
DRAM[21624] = 8'b10111110;
DRAM[21625] = 8'b10110101;
DRAM[21626] = 8'b10111110;
DRAM[21627] = 8'b10110011;
DRAM[21628] = 8'b10111000;
DRAM[21629] = 8'b10111110;
DRAM[21630] = 8'b10101101;
DRAM[21631] = 8'b11000010;
DRAM[21632] = 8'b10110101;
DRAM[21633] = 8'b10101100;
DRAM[21634] = 8'b10101110;
DRAM[21635] = 8'b10111110;
DRAM[21636] = 8'b11001000;
DRAM[21637] = 8'b11001011;
DRAM[21638] = 8'b11000010;
DRAM[21639] = 8'b10101000;
DRAM[21640] = 8'b11000000;
DRAM[21641] = 8'b11001111;
DRAM[21642] = 8'b10111100;
DRAM[21643] = 8'b10110000;
DRAM[21644] = 8'b11000101;
DRAM[21645] = 8'b11000111;
DRAM[21646] = 8'b10110110;
DRAM[21647] = 8'b10111010;
DRAM[21648] = 8'b10110100;
DRAM[21649] = 8'b10111010;
DRAM[21650] = 8'b10110110;
DRAM[21651] = 8'b10110000;
DRAM[21652] = 8'b10101100;
DRAM[21653] = 8'b10100010;
DRAM[21654] = 8'b10100011;
DRAM[21655] = 8'b10110001;
DRAM[21656] = 8'b10101101;
DRAM[21657] = 8'b10111110;
DRAM[21658] = 8'b10101110;
DRAM[21659] = 8'b10100010;
DRAM[21660] = 8'b10110110;
DRAM[21661] = 8'b10110101;
DRAM[21662] = 8'b10100100;
DRAM[21663] = 8'b10100111;
DRAM[21664] = 8'b11001100;
DRAM[21665] = 8'b11001100;
DRAM[21666] = 8'b10111101;
DRAM[21667] = 8'b10110101;
DRAM[21668] = 8'b10111110;
DRAM[21669] = 8'b11000100;
DRAM[21670] = 8'b11000001;
DRAM[21671] = 8'b11000010;
DRAM[21672] = 8'b11000101;
DRAM[21673] = 8'b11001100;
DRAM[21674] = 8'b11010100;
DRAM[21675] = 8'b11010101;
DRAM[21676] = 8'b11001110;
DRAM[21677] = 8'b11000100;
DRAM[21678] = 8'b10111110;
DRAM[21679] = 8'b10111011;
DRAM[21680] = 8'b11000110;
DRAM[21681] = 8'b11001010;
DRAM[21682] = 8'b11010000;
DRAM[21683] = 8'b11010110;
DRAM[21684] = 8'b11011011;
DRAM[21685] = 8'b11011111;
DRAM[21686] = 8'b11100010;
DRAM[21687] = 8'b11100100;
DRAM[21688] = 8'b11010000;
DRAM[21689] = 8'b11010111;
DRAM[21690] = 8'b11010111;
DRAM[21691] = 8'b11001111;
DRAM[21692] = 8'b11001100;
DRAM[21693] = 8'b11000101;
DRAM[21694] = 8'b10101110;
DRAM[21695] = 8'b10010011;
DRAM[21696] = 8'b1110011;
DRAM[21697] = 8'b1101011;
DRAM[21698] = 8'b1000010;
DRAM[21699] = 8'b1101111;
DRAM[21700] = 8'b10000111;
DRAM[21701] = 8'b10100000;
DRAM[21702] = 8'b10010010;
DRAM[21703] = 8'b11000111;
DRAM[21704] = 8'b10110100;
DRAM[21705] = 8'b11010111;
DRAM[21706] = 8'b11101111;
DRAM[21707] = 8'b11111001;
DRAM[21708] = 8'b11111111;
DRAM[21709] = 8'b11110101;
DRAM[21710] = 8'b11101010;
DRAM[21711] = 8'b11101111;
DRAM[21712] = 8'b11100011;
DRAM[21713] = 8'b11000000;
DRAM[21714] = 8'b11001110;
DRAM[21715] = 8'b11100011;
DRAM[21716] = 8'b11001110;
DRAM[21717] = 8'b11000100;
DRAM[21718] = 8'b11001110;
DRAM[21719] = 8'b11010110;
DRAM[21720] = 8'b11010101;
DRAM[21721] = 8'b11001000;
DRAM[21722] = 8'b11001000;
DRAM[21723] = 8'b10111101;
DRAM[21724] = 8'b11101010;
DRAM[21725] = 8'b11010111;
DRAM[21726] = 8'b11000111;
DRAM[21727] = 8'b11100100;
DRAM[21728] = 8'b11011111;
DRAM[21729] = 8'b11100111;
DRAM[21730] = 8'b11101110;
DRAM[21731] = 8'b11100010;
DRAM[21732] = 8'b11011101;
DRAM[21733] = 8'b11110111;
DRAM[21734] = 8'b11111111;
DRAM[21735] = 8'b11100101;
DRAM[21736] = 8'b11110010;
DRAM[21737] = 8'b11110110;
DRAM[21738] = 8'b10110111;
DRAM[21739] = 8'b10100011;
DRAM[21740] = 8'b10000010;
DRAM[21741] = 8'b1110010;
DRAM[21742] = 8'b1101101;
DRAM[21743] = 8'b1101110;
DRAM[21744] = 8'b1101001;
DRAM[21745] = 8'b1100111;
DRAM[21746] = 8'b1100101;
DRAM[21747] = 8'b1100101;
DRAM[21748] = 8'b1100110;
DRAM[21749] = 8'b1100110;
DRAM[21750] = 8'b1100100;
DRAM[21751] = 8'b1100010;
DRAM[21752] = 8'b1100011;
DRAM[21753] = 8'b1100011;
DRAM[21754] = 8'b1100010;
DRAM[21755] = 8'b1100010;
DRAM[21756] = 8'b1100001;
DRAM[21757] = 8'b1100001;
DRAM[21758] = 8'b1100000;
DRAM[21759] = 8'b1100000;
DRAM[21760] = 8'b1110101;
DRAM[21761] = 8'b1110101;
DRAM[21762] = 8'b1110110;
DRAM[21763] = 8'b1110110;
DRAM[21764] = 8'b1110110;
DRAM[21765] = 8'b1110111;
DRAM[21766] = 8'b1110111;
DRAM[21767] = 8'b1110111;
DRAM[21768] = 8'b1111001;
DRAM[21769] = 8'b1111001;
DRAM[21770] = 8'b1111010;
DRAM[21771] = 8'b1111010;
DRAM[21772] = 8'b1111010;
DRAM[21773] = 8'b1111011;
DRAM[21774] = 8'b1111011;
DRAM[21775] = 8'b1111011;
DRAM[21776] = 8'b1111111;
DRAM[21777] = 8'b1111101;
DRAM[21778] = 8'b1111010;
DRAM[21779] = 8'b1111000;
DRAM[21780] = 8'b1111011;
DRAM[21781] = 8'b10000100;
DRAM[21782] = 8'b10010000;
DRAM[21783] = 8'b10011001;
DRAM[21784] = 8'b10011111;
DRAM[21785] = 8'b10111000;
DRAM[21786] = 8'b11011000;
DRAM[21787] = 8'b11101111;
DRAM[21788] = 8'b11111011;
DRAM[21789] = 8'b11111111;
DRAM[21790] = 8'b11111101;
DRAM[21791] = 8'b11111000;
DRAM[21792] = 8'b11111111;
DRAM[21793] = 8'b11111001;
DRAM[21794] = 8'b11110010;
DRAM[21795] = 8'b11110000;
DRAM[21796] = 8'b11110011;
DRAM[21797] = 8'b11110110;
DRAM[21798] = 8'b11110101;
DRAM[21799] = 8'b11110011;
DRAM[21800] = 8'b11100110;
DRAM[21801] = 8'b11101000;
DRAM[21802] = 8'b11100100;
DRAM[21803] = 8'b11011100;
DRAM[21804] = 8'b11011010;
DRAM[21805] = 8'b11011111;
DRAM[21806] = 8'b11100110;
DRAM[21807] = 8'b11101010;
DRAM[21808] = 8'b11100100;
DRAM[21809] = 8'b11011000;
DRAM[21810] = 8'b11101101;
DRAM[21811] = 8'b11100100;
DRAM[21812] = 8'b11100110;
DRAM[21813] = 8'b11110001;
DRAM[21814] = 8'b11011001;
DRAM[21815] = 8'b11100001;
DRAM[21816] = 8'b11100000;
DRAM[21817] = 8'b11011101;
DRAM[21818] = 8'b11010110;
DRAM[21819] = 8'b11100000;
DRAM[21820] = 8'b11101000;
DRAM[21821] = 8'b11010100;
DRAM[21822] = 8'b11010000;
DRAM[21823] = 8'b11101110;
DRAM[21824] = 8'b11100000;
DRAM[21825] = 8'b11100110;
DRAM[21826] = 8'b11110110;
DRAM[21827] = 8'b11100111;
DRAM[21828] = 8'b11100110;
DRAM[21829] = 8'b11110101;
DRAM[21830] = 8'b11100110;
DRAM[21831] = 8'b11010000;
DRAM[21832] = 8'b11000101;
DRAM[21833] = 8'b10111110;
DRAM[21834] = 8'b10101001;
DRAM[21835] = 8'b10101011;
DRAM[21836] = 8'b10001100;
DRAM[21837] = 8'b1011110;
DRAM[21838] = 8'b1000101;
DRAM[21839] = 8'b1100111;
DRAM[21840] = 8'b1101000;
DRAM[21841] = 8'b1110111;
DRAM[21842] = 8'b10001010;
DRAM[21843] = 8'b10010101;
DRAM[21844] = 8'b10011011;
DRAM[21845] = 8'b10100100;
DRAM[21846] = 8'b10110011;
DRAM[21847] = 8'b11000000;
DRAM[21848] = 8'b11001110;
DRAM[21849] = 8'b11010000;
DRAM[21850] = 8'b11010011;
DRAM[21851] = 8'b11010101;
DRAM[21852] = 8'b11010110;
DRAM[21853] = 8'b11011000;
DRAM[21854] = 8'b11011010;
DRAM[21855] = 8'b11011100;
DRAM[21856] = 8'b11011111;
DRAM[21857] = 8'b11001111;
DRAM[21858] = 8'b11000100;
DRAM[21859] = 8'b11001000;
DRAM[21860] = 8'b11010101;
DRAM[21861] = 8'b11010101;
DRAM[21862] = 8'b11000010;
DRAM[21863] = 8'b10101110;
DRAM[21864] = 8'b10111001;
DRAM[21865] = 8'b10111000;
DRAM[21866] = 8'b10111100;
DRAM[21867] = 8'b11000110;
DRAM[21868] = 8'b11001101;
DRAM[21869] = 8'b11001010;
DRAM[21870] = 8'b10111011;
DRAM[21871] = 8'b10101110;
DRAM[21872] = 8'b10110100;
DRAM[21873] = 8'b10111001;
DRAM[21874] = 8'b10111100;
DRAM[21875] = 8'b10111010;
DRAM[21876] = 8'b10110011;
DRAM[21877] = 8'b10101110;
DRAM[21878] = 8'b10101101;
DRAM[21879] = 8'b10101110;
DRAM[21880] = 8'b10110100;
DRAM[21881] = 8'b10101110;
DRAM[21882] = 8'b10101111;
DRAM[21883] = 8'b10110000;
DRAM[21884] = 8'b10111101;
DRAM[21885] = 8'b11000000;
DRAM[21886] = 8'b10110101;
DRAM[21887] = 8'b11000000;
DRAM[21888] = 8'b10111000;
DRAM[21889] = 8'b10101110;
DRAM[21890] = 8'b10100011;
DRAM[21891] = 8'b10110100;
DRAM[21892] = 8'b11000011;
DRAM[21893] = 8'b11001000;
DRAM[21894] = 8'b11000100;
DRAM[21895] = 8'b10100100;
DRAM[21896] = 8'b10111010;
DRAM[21897] = 8'b11000000;
DRAM[21898] = 8'b10110001;
DRAM[21899] = 8'b10101010;
DRAM[21900] = 8'b10111101;
DRAM[21901] = 8'b11000100;
DRAM[21902] = 8'b10111000;
DRAM[21903] = 8'b10110100;
DRAM[21904] = 8'b10110000;
DRAM[21905] = 8'b10110100;
DRAM[21906] = 8'b10101110;
DRAM[21907] = 8'b10101010;
DRAM[21908] = 8'b10101010;
DRAM[21909] = 8'b10100100;
DRAM[21910] = 8'b10100100;
DRAM[21911] = 8'b10110001;
DRAM[21912] = 8'b10101001;
DRAM[21913] = 8'b10110101;
DRAM[21914] = 8'b10101000;
DRAM[21915] = 8'b10011010;
DRAM[21916] = 8'b10100110;
DRAM[21917] = 8'b10101101;
DRAM[21918] = 8'b10101110;
DRAM[21919] = 8'b10111000;
DRAM[21920] = 8'b11000101;
DRAM[21921] = 8'b11000011;
DRAM[21922] = 8'b10110101;
DRAM[21923] = 8'b10110001;
DRAM[21924] = 8'b11000001;
DRAM[21925] = 8'b11001001;
DRAM[21926] = 8'b11000101;
DRAM[21927] = 8'b11000011;
DRAM[21928] = 8'b11010000;
DRAM[21929] = 8'b11001101;
DRAM[21930] = 8'b11000101;
DRAM[21931] = 8'b10111010;
DRAM[21932] = 8'b10110011;
DRAM[21933] = 8'b10111000;
DRAM[21934] = 8'b11000111;
DRAM[21935] = 8'b11010011;
DRAM[21936] = 8'b11000111;
DRAM[21937] = 8'b11001000;
DRAM[21938] = 8'b11001011;
DRAM[21939] = 8'b11010000;
DRAM[21940] = 8'b11010100;
DRAM[21941] = 8'b11010100;
DRAM[21942] = 8'b11010010;
DRAM[21943] = 8'b11001111;
DRAM[21944] = 8'b11011000;
DRAM[21945] = 8'b11010110;
DRAM[21946] = 8'b11010011;
DRAM[21947] = 8'b11010000;
DRAM[21948] = 8'b11001111;
DRAM[21949] = 8'b11000111;
DRAM[21950] = 8'b10110100;
DRAM[21951] = 8'b10100010;
DRAM[21952] = 8'b10000111;
DRAM[21953] = 8'b1101001;
DRAM[21954] = 8'b110011;
DRAM[21955] = 8'b1101011;
DRAM[21956] = 8'b10000000;
DRAM[21957] = 8'b10011001;
DRAM[21958] = 8'b10001111;
DRAM[21959] = 8'b11010000;
DRAM[21960] = 8'b10110101;
DRAM[21961] = 8'b11001000;
DRAM[21962] = 8'b11100110;
DRAM[21963] = 8'b11111011;
DRAM[21964] = 8'b11111100;
DRAM[21965] = 8'b11110110;
DRAM[21966] = 8'b11101110;
DRAM[21967] = 8'b11100110;
DRAM[21968] = 8'b11111011;
DRAM[21969] = 8'b10111110;
DRAM[21970] = 8'b11001010;
DRAM[21971] = 8'b11001100;
DRAM[21972] = 8'b11100010;
DRAM[21973] = 8'b11001100;
DRAM[21974] = 8'b11001101;
DRAM[21975] = 8'b11000101;
DRAM[21976] = 8'b11010011;
DRAM[21977] = 8'b11000010;
DRAM[21978] = 8'b10111010;
DRAM[21979] = 8'b11000010;
DRAM[21980] = 8'b11001100;
DRAM[21981] = 8'b11100000;
DRAM[21982] = 8'b10111001;
DRAM[21983] = 8'b11010111;
DRAM[21984] = 8'b11100010;
DRAM[21985] = 8'b11010110;
DRAM[21986] = 8'b11100111;
DRAM[21987] = 8'b11101011;
DRAM[21988] = 8'b11010001;
DRAM[21989] = 8'b11010110;
DRAM[21990] = 8'b11110010;
DRAM[21991] = 8'b11110011;
DRAM[21992] = 8'b11111001;
DRAM[21993] = 8'b11111010;
DRAM[21994] = 8'b11000110;
DRAM[21995] = 8'b10100011;
DRAM[21996] = 8'b10001101;
DRAM[21997] = 8'b1111001;
DRAM[21998] = 8'b1101000;
DRAM[21999] = 8'b1101001;
DRAM[22000] = 8'b1101001;
DRAM[22001] = 8'b1101000;
DRAM[22002] = 8'b1100110;
DRAM[22003] = 8'b1100110;
DRAM[22004] = 8'b1100111;
DRAM[22005] = 8'b1100110;
DRAM[22006] = 8'b1100101;
DRAM[22007] = 8'b1100011;
DRAM[22008] = 8'b1100100;
DRAM[22009] = 8'b1100100;
DRAM[22010] = 8'b1100011;
DRAM[22011] = 8'b1100011;
DRAM[22012] = 8'b1100010;
DRAM[22013] = 8'b1100001;
DRAM[22014] = 8'b1100001;
DRAM[22015] = 8'b1100000;
DRAM[22016] = 8'b1110111;
DRAM[22017] = 8'b1110111;
DRAM[22018] = 8'b1111000;
DRAM[22019] = 8'b1111000;
DRAM[22020] = 8'b1111000;
DRAM[22021] = 8'b1111001;
DRAM[22022] = 8'b1111001;
DRAM[22023] = 8'b1111001;
DRAM[22024] = 8'b1111010;
DRAM[22025] = 8'b1111010;
DRAM[22026] = 8'b1111010;
DRAM[22027] = 8'b1111011;
DRAM[22028] = 8'b1111011;
DRAM[22029] = 8'b1111011;
DRAM[22030] = 8'b1111100;
DRAM[22031] = 8'b1111100;
DRAM[22032] = 8'b1111110;
DRAM[22033] = 8'b1111101;
DRAM[22034] = 8'b1111011;
DRAM[22035] = 8'b1111010;
DRAM[22036] = 8'b1111100;
DRAM[22037] = 8'b10000101;
DRAM[22038] = 8'b10001111;
DRAM[22039] = 8'b10010111;
DRAM[22040] = 8'b10011000;
DRAM[22041] = 8'b11001000;
DRAM[22042] = 8'b11110000;
DRAM[22043] = 8'b11110101;
DRAM[22044] = 8'b11110010;
DRAM[22045] = 8'b11111001;
DRAM[22046] = 8'b11111100;
DRAM[22047] = 8'b11110110;
DRAM[22048] = 8'b11111001;
DRAM[22049] = 8'b11110011;
DRAM[22050] = 8'b11101110;
DRAM[22051] = 8'b11101111;
DRAM[22052] = 8'b11110011;
DRAM[22053] = 8'b11110101;
DRAM[22054] = 8'b11110001;
DRAM[22055] = 8'b11101011;
DRAM[22056] = 8'b11011111;
DRAM[22057] = 8'b11101000;
DRAM[22058] = 8'b11100111;
DRAM[22059] = 8'b11011110;
DRAM[22060] = 8'b11011101;
DRAM[22061] = 8'b11100110;
DRAM[22062] = 8'b11100100;
DRAM[22063] = 8'b11011000;
DRAM[22064] = 8'b11010101;
DRAM[22065] = 8'b11011101;
DRAM[22066] = 8'b11101001;
DRAM[22067] = 8'b11100111;
DRAM[22068] = 8'b11100010;
DRAM[22069] = 8'b11100011;
DRAM[22070] = 8'b11100010;
DRAM[22071] = 8'b11101000;
DRAM[22072] = 8'b11011001;
DRAM[22073] = 8'b11010001;
DRAM[22074] = 8'b11011101;
DRAM[22075] = 8'b11101010;
DRAM[22076] = 8'b11011101;
DRAM[22077] = 8'b11010000;
DRAM[22078] = 8'b11011001;
DRAM[22079] = 8'b11100101;
DRAM[22080] = 8'b11011011;
DRAM[22081] = 8'b11101011;
DRAM[22082] = 8'b11101110;
DRAM[22083] = 8'b11100100;
DRAM[22084] = 8'b11100010;
DRAM[22085] = 8'b11111110;
DRAM[22086] = 8'b11011100;
DRAM[22087] = 8'b11010011;
DRAM[22088] = 8'b11010010;
DRAM[22089] = 8'b10110111;
DRAM[22090] = 8'b10101011;
DRAM[22091] = 8'b10011111;
DRAM[22092] = 8'b10000111;
DRAM[22093] = 8'b1010100;
DRAM[22094] = 8'b1001101;
DRAM[22095] = 8'b1011110;
DRAM[22096] = 8'b1111000;
DRAM[22097] = 8'b10001010;
DRAM[22098] = 8'b10100100;
DRAM[22099] = 8'b10111000;
DRAM[22100] = 8'b11000100;
DRAM[22101] = 8'b11001011;
DRAM[22102] = 8'b11010011;
DRAM[22103] = 8'b11011000;
DRAM[22104] = 8'b11000110;
DRAM[22105] = 8'b11010101;
DRAM[22106] = 8'b11100101;
DRAM[22107] = 8'b11101000;
DRAM[22108] = 8'b11011111;
DRAM[22109] = 8'b11010110;
DRAM[22110] = 8'b11010110;
DRAM[22111] = 8'b11011010;
DRAM[22112] = 8'b11010101;
DRAM[22113] = 8'b11100011;
DRAM[22114] = 8'b11101010;
DRAM[22115] = 8'b11011100;
DRAM[22116] = 8'b11000110;
DRAM[22117] = 8'b10111111;
DRAM[22118] = 8'b11010001;
DRAM[22119] = 8'b11100110;
DRAM[22120] = 8'b10111110;
DRAM[22121] = 8'b10110110;
DRAM[22122] = 8'b10110010;
DRAM[22123] = 8'b10111010;
DRAM[22124] = 8'b11000111;
DRAM[22125] = 8'b11001101;
DRAM[22126] = 8'b11000101;
DRAM[22127] = 8'b10111011;
DRAM[22128] = 8'b10111000;
DRAM[22129] = 8'b10111101;
DRAM[22130] = 8'b10111011;
DRAM[22131] = 8'b10110100;
DRAM[22132] = 8'b10110000;
DRAM[22133] = 8'b10110001;
DRAM[22134] = 8'b10101011;
DRAM[22135] = 8'b10100001;
DRAM[22136] = 8'b10101100;
DRAM[22137] = 8'b10110011;
DRAM[22138] = 8'b10100110;
DRAM[22139] = 8'b10101100;
DRAM[22140] = 8'b11000010;
DRAM[22141] = 8'b11000111;
DRAM[22142] = 8'b10111110;
DRAM[22143] = 8'b10101100;
DRAM[22144] = 8'b10111000;
DRAM[22145] = 8'b10110001;
DRAM[22146] = 8'b10011111;
DRAM[22147] = 8'b10101101;
DRAM[22148] = 8'b10110111;
DRAM[22149] = 8'b10111100;
DRAM[22150] = 8'b11000010;
DRAM[22151] = 8'b10100100;
DRAM[22152] = 8'b10110111;
DRAM[22153] = 8'b10111000;
DRAM[22154] = 8'b10110001;
DRAM[22155] = 8'b10101100;
DRAM[22156] = 8'b10110100;
DRAM[22157] = 8'b10111110;
DRAM[22158] = 8'b10111011;
DRAM[22159] = 8'b10110001;
DRAM[22160] = 8'b10101100;
DRAM[22161] = 8'b10101101;
DRAM[22162] = 8'b10101000;
DRAM[22163] = 8'b10100111;
DRAM[22164] = 8'b10101100;
DRAM[22165] = 8'b10100101;
DRAM[22166] = 8'b10100000;
DRAM[22167] = 8'b10101000;
DRAM[22168] = 8'b10100001;
DRAM[22169] = 8'b10101011;
DRAM[22170] = 8'b10101011;
DRAM[22171] = 8'b10100000;
DRAM[22172] = 8'b10011110;
DRAM[22173] = 8'b10101001;
DRAM[22174] = 8'b10110111;
DRAM[22175] = 8'b11000000;
DRAM[22176] = 8'b10101101;
DRAM[22177] = 8'b10101110;
DRAM[22178] = 8'b10100101;
DRAM[22179] = 8'b10100110;
DRAM[22180] = 8'b10111010;
DRAM[22181] = 8'b11000111;
DRAM[22182] = 8'b11000111;
DRAM[22183] = 8'b11001001;
DRAM[22184] = 8'b10110110;
DRAM[22185] = 8'b10111101;
DRAM[22186] = 8'b11000111;
DRAM[22187] = 8'b11001110;
DRAM[22188] = 8'b11010000;
DRAM[22189] = 8'b11010000;
DRAM[22190] = 8'b11010000;
DRAM[22191] = 8'b11010001;
DRAM[22192] = 8'b11001001;
DRAM[22193] = 8'b11000110;
DRAM[22194] = 8'b11000101;
DRAM[22195] = 8'b11001010;
DRAM[22196] = 8'b11010000;
DRAM[22197] = 8'b11010010;
DRAM[22198] = 8'b11001110;
DRAM[22199] = 8'b11001000;
DRAM[22200] = 8'b11010101;
DRAM[22201] = 8'b11010000;
DRAM[22202] = 8'b11001101;
DRAM[22203] = 8'b11001100;
DRAM[22204] = 8'b11000010;
DRAM[22205] = 8'b10101101;
DRAM[22206] = 8'b10011000;
DRAM[22207] = 8'b10001101;
DRAM[22208] = 8'b1101111;
DRAM[22209] = 8'b1010101;
DRAM[22210] = 8'b111011;
DRAM[22211] = 8'b1100110;
DRAM[22212] = 8'b10001100;
DRAM[22213] = 8'b10010111;
DRAM[22214] = 8'b10001111;
DRAM[22215] = 8'b10101101;
DRAM[22216] = 8'b10111101;
DRAM[22217] = 8'b11000001;
DRAM[22218] = 8'b11100101;
DRAM[22219] = 8'b11111111;
DRAM[22220] = 8'b11111000;
DRAM[22221] = 8'b11111001;
DRAM[22222] = 8'b11111100;
DRAM[22223] = 8'b11101010;
DRAM[22224] = 8'b11111001;
DRAM[22225] = 8'b11000111;
DRAM[22226] = 8'b11000111;
DRAM[22227] = 8'b11001000;
DRAM[22228] = 8'b11011011;
DRAM[22229] = 8'b11010000;
DRAM[22230] = 8'b11000100;
DRAM[22231] = 8'b11001110;
DRAM[22232] = 8'b11010010;
DRAM[22233] = 8'b10111100;
DRAM[22234] = 8'b10110011;
DRAM[22235] = 8'b11000110;
DRAM[22236] = 8'b10110111;
DRAM[22237] = 8'b11010001;
DRAM[22238] = 8'b11001110;
DRAM[22239] = 8'b11001101;
DRAM[22240] = 8'b11011010;
DRAM[22241] = 8'b11010010;
DRAM[22242] = 8'b11010110;
DRAM[22243] = 8'b11011010;
DRAM[22244] = 8'b11010010;
DRAM[22245] = 8'b11010000;
DRAM[22246] = 8'b11100010;
DRAM[22247] = 8'b11110100;
DRAM[22248] = 8'b11111010;
DRAM[22249] = 8'b11111010;
DRAM[22250] = 8'b11011011;
DRAM[22251] = 8'b10100000;
DRAM[22252] = 8'b10010100;
DRAM[22253] = 8'b1111110;
DRAM[22254] = 8'b1100110;
DRAM[22255] = 8'b1101100;
DRAM[22256] = 8'b1101010;
DRAM[22257] = 8'b1101000;
DRAM[22258] = 8'b1100111;
DRAM[22259] = 8'b1100110;
DRAM[22260] = 8'b1100111;
DRAM[22261] = 8'b1100111;
DRAM[22262] = 8'b1100101;
DRAM[22263] = 8'b1100011;
DRAM[22264] = 8'b1100101;
DRAM[22265] = 8'b1100101;
DRAM[22266] = 8'b1100100;
DRAM[22267] = 8'b1100011;
DRAM[22268] = 8'b1100010;
DRAM[22269] = 8'b1100001;
DRAM[22270] = 8'b1100001;
DRAM[22271] = 8'b1100000;
DRAM[22272] = 8'b1111000;
DRAM[22273] = 8'b1111000;
DRAM[22274] = 8'b1111001;
DRAM[22275] = 8'b1111001;
DRAM[22276] = 8'b1111001;
DRAM[22277] = 8'b1111010;
DRAM[22278] = 8'b1111010;
DRAM[22279] = 8'b1111010;
DRAM[22280] = 8'b1111010;
DRAM[22281] = 8'b1111010;
DRAM[22282] = 8'b1111011;
DRAM[22283] = 8'b1111011;
DRAM[22284] = 8'b1111011;
DRAM[22285] = 8'b1111100;
DRAM[22286] = 8'b1111100;
DRAM[22287] = 8'b1111100;
DRAM[22288] = 8'b1111001;
DRAM[22289] = 8'b1111011;
DRAM[22290] = 8'b1111110;
DRAM[22291] = 8'b10000000;
DRAM[22292] = 8'b10000001;
DRAM[22293] = 8'b10000010;
DRAM[22294] = 8'b10000100;
DRAM[22295] = 8'b10000111;
DRAM[22296] = 8'b10100111;
DRAM[22297] = 8'b10101100;
DRAM[22298] = 8'b11001011;
DRAM[22299] = 8'b11110010;
DRAM[22300] = 8'b11111011;
DRAM[22301] = 8'b11101010;
DRAM[22302] = 8'b11101001;
DRAM[22303] = 8'b11111011;
DRAM[22304] = 8'b11110011;
DRAM[22305] = 8'b11101111;
DRAM[22306] = 8'b11101101;
DRAM[22307] = 8'b11110000;
DRAM[22308] = 8'b11110101;
DRAM[22309] = 8'b11110101;
DRAM[22310] = 8'b11101101;
DRAM[22311] = 8'b11100110;
DRAM[22312] = 8'b11011111;
DRAM[22313] = 8'b11101101;
DRAM[22314] = 8'b11101110;
DRAM[22315] = 8'b11100011;
DRAM[22316] = 8'b11100100;
DRAM[22317] = 8'b11101010;
DRAM[22318] = 8'b11011011;
DRAM[22319] = 8'b11000001;
DRAM[22320] = 8'b11010101;
DRAM[22321] = 8'b11101101;
DRAM[22322] = 8'b11011010;
DRAM[22323] = 8'b11010110;
DRAM[22324] = 8'b11011101;
DRAM[22325] = 8'b11100100;
DRAM[22326] = 8'b11101000;
DRAM[22327] = 8'b11000000;
DRAM[22328] = 8'b11010010;
DRAM[22329] = 8'b11001101;
DRAM[22330] = 8'b11101000;
DRAM[22331] = 8'b11101000;
DRAM[22332] = 8'b11001001;
DRAM[22333] = 8'b11011010;
DRAM[22334] = 8'b11101011;
DRAM[22335] = 8'b11000110;
DRAM[22336] = 8'b11011111;
DRAM[22337] = 8'b11101101;
DRAM[22338] = 8'b11110100;
DRAM[22339] = 8'b11011011;
DRAM[22340] = 8'b11101101;
DRAM[22341] = 8'b11111110;
DRAM[22342] = 8'b11011010;
DRAM[22343] = 8'b11010000;
DRAM[22344] = 8'b11011011;
DRAM[22345] = 8'b10110011;
DRAM[22346] = 8'b10101101;
DRAM[22347] = 8'b10011011;
DRAM[22348] = 8'b10001101;
DRAM[22349] = 8'b1011101;
DRAM[22350] = 8'b1100011;
DRAM[22351] = 8'b1101000;
DRAM[22352] = 8'b1100010;
DRAM[22353] = 8'b1101110;
DRAM[22354] = 8'b10000001;
DRAM[22355] = 8'b10010111;
DRAM[22356] = 8'b10101100;
DRAM[22357] = 8'b10111110;
DRAM[22358] = 8'b11001100;
DRAM[22359] = 8'b11010011;
DRAM[22360] = 8'b11100100;
DRAM[22361] = 8'b11011111;
DRAM[22362] = 8'b11011100;
DRAM[22363] = 8'b11100000;
DRAM[22364] = 8'b11100110;
DRAM[22365] = 8'b11100111;
DRAM[22366] = 8'b11100000;
DRAM[22367] = 8'b11011000;
DRAM[22368] = 8'b11001111;
DRAM[22369] = 8'b11000111;
DRAM[22370] = 8'b10111111;
DRAM[22371] = 8'b10111110;
DRAM[22372] = 8'b11000011;
DRAM[22373] = 8'b11001001;
DRAM[22374] = 8'b11001010;
DRAM[22375] = 8'b11001000;
DRAM[22376] = 8'b11010111;
DRAM[22377] = 8'b11001100;
DRAM[22378] = 8'b10111110;
DRAM[22379] = 8'b10110100;
DRAM[22380] = 8'b10110011;
DRAM[22381] = 8'b10111001;
DRAM[22382] = 8'b11000001;
DRAM[22383] = 8'b11000110;
DRAM[22384] = 8'b10111000;
DRAM[22385] = 8'b10111110;
DRAM[22386] = 8'b10111011;
DRAM[22387] = 8'b10110100;
DRAM[22388] = 8'b10111000;
DRAM[22389] = 8'b11000010;
DRAM[22390] = 8'b10111101;
DRAM[22391] = 8'b10101110;
DRAM[22392] = 8'b10011010;
DRAM[22393] = 8'b11000010;
DRAM[22394] = 8'b10111001;
DRAM[22395] = 8'b10110110;
DRAM[22396] = 8'b10111011;
DRAM[22397] = 8'b10111010;
DRAM[22398] = 8'b11000000;
DRAM[22399] = 8'b10101000;
DRAM[22400] = 8'b10110111;
DRAM[22401] = 8'b10110100;
DRAM[22402] = 8'b10011111;
DRAM[22403] = 8'b10101000;
DRAM[22404] = 8'b10101101;
DRAM[22405] = 8'b10110001;
DRAM[22406] = 8'b10111111;
DRAM[22407] = 8'b10100100;
DRAM[22408] = 8'b10111010;
DRAM[22409] = 8'b10111000;
DRAM[22410] = 8'b10110111;
DRAM[22411] = 8'b10110010;
DRAM[22412] = 8'b10101110;
DRAM[22413] = 8'b10111000;
DRAM[22414] = 8'b10111100;
DRAM[22415] = 8'b10110000;
DRAM[22416] = 8'b10101001;
DRAM[22417] = 8'b10101010;
DRAM[22418] = 8'b10100100;
DRAM[22419] = 8'b10100110;
DRAM[22420] = 8'b10101110;
DRAM[22421] = 8'b10100110;
DRAM[22422] = 8'b10011100;
DRAM[22423] = 8'b10011111;
DRAM[22424] = 8'b10010101;
DRAM[22425] = 8'b10100010;
DRAM[22426] = 8'b10110001;
DRAM[22427] = 8'b10101100;
DRAM[22428] = 8'b10100001;
DRAM[22429] = 8'b10101010;
DRAM[22430] = 8'b10111010;
DRAM[22431] = 8'b10111101;
DRAM[22432] = 8'b10101011;
DRAM[22433] = 8'b10101110;
DRAM[22434] = 8'b10100100;
DRAM[22435] = 8'b10011111;
DRAM[22436] = 8'b10101011;
DRAM[22437] = 8'b10110100;
DRAM[22438] = 8'b10110101;
DRAM[22439] = 8'b10111001;
DRAM[22440] = 8'b11000001;
DRAM[22441] = 8'b11000101;
DRAM[22442] = 8'b11001101;
DRAM[22443] = 8'b11010100;
DRAM[22444] = 8'b11011000;
DRAM[22445] = 8'b11010101;
DRAM[22446] = 8'b11001110;
DRAM[22447] = 8'b11001000;
DRAM[22448] = 8'b11001001;
DRAM[22449] = 8'b11000100;
DRAM[22450] = 8'b11000010;
DRAM[22451] = 8'b11001001;
DRAM[22452] = 8'b11010100;
DRAM[22453] = 8'b11011011;
DRAM[22454] = 8'b11011000;
DRAM[22455] = 8'b11010010;
DRAM[22456] = 8'b11011001;
DRAM[22457] = 8'b11010111;
DRAM[22458] = 8'b11011100;
DRAM[22459] = 8'b11011111;
DRAM[22460] = 8'b11001101;
DRAM[22461] = 8'b10101010;
DRAM[22462] = 8'b10010000;
DRAM[22463] = 8'b10001001;
DRAM[22464] = 8'b1111001;
DRAM[22465] = 8'b1011111;
DRAM[22466] = 8'b1001001;
DRAM[22467] = 8'b1000001;
DRAM[22468] = 8'b1111000;
DRAM[22469] = 8'b10001111;
DRAM[22470] = 8'b10100000;
DRAM[22471] = 8'b10011101;
DRAM[22472] = 8'b11000001;
DRAM[22473] = 8'b10111011;
DRAM[22474] = 8'b11100011;
DRAM[22475] = 8'b11111111;
DRAM[22476] = 8'b11110000;
DRAM[22477] = 8'b11110111;
DRAM[22478] = 8'b11111111;
DRAM[22479] = 8'b11101110;
DRAM[22480] = 8'b11100110;
DRAM[22481] = 8'b11010110;
DRAM[22482] = 8'b11000100;
DRAM[22483] = 8'b11011000;
DRAM[22484] = 8'b10111111;
DRAM[22485] = 8'b11010010;
DRAM[22486] = 8'b10110101;
DRAM[22487] = 8'b11100100;
DRAM[22488] = 8'b11001001;
DRAM[22489] = 8'b11011011;
DRAM[22490] = 8'b10110111;
DRAM[22491] = 8'b10100111;
DRAM[22492] = 8'b11010000;
DRAM[22493] = 8'b10111000;
DRAM[22494] = 8'b11000111;
DRAM[22495] = 8'b11010000;
DRAM[22496] = 8'b11001110;
DRAM[22497] = 8'b11010111;
DRAM[22498] = 8'b11000100;
DRAM[22499] = 8'b10111100;
DRAM[22500] = 8'b11011000;
DRAM[22501] = 8'b11100100;
DRAM[22502] = 8'b11011110;
DRAM[22503] = 8'b11101000;
DRAM[22504] = 8'b11110001;
DRAM[22505] = 8'b11110001;
DRAM[22506] = 8'b11100011;
DRAM[22507] = 8'b10010111;
DRAM[22508] = 8'b10010001;
DRAM[22509] = 8'b1111100;
DRAM[22510] = 8'b1100010;
DRAM[22511] = 8'b1101110;
DRAM[22512] = 8'b1101010;
DRAM[22513] = 8'b1101001;
DRAM[22514] = 8'b1100111;
DRAM[22515] = 8'b1100111;
DRAM[22516] = 8'b1100111;
DRAM[22517] = 8'b1100111;
DRAM[22518] = 8'b1100110;
DRAM[22519] = 8'b1100100;
DRAM[22520] = 8'b1100110;
DRAM[22521] = 8'b1100101;
DRAM[22522] = 8'b1100100;
DRAM[22523] = 8'b1100100;
DRAM[22524] = 8'b1100011;
DRAM[22525] = 8'b1100010;
DRAM[22526] = 8'b1100001;
DRAM[22527] = 8'b1100001;
DRAM[22528] = 8'b1111001;
DRAM[22529] = 8'b1111001;
DRAM[22530] = 8'b1111001;
DRAM[22531] = 8'b1111010;
DRAM[22532] = 8'b1111010;
DRAM[22533] = 8'b1111011;
DRAM[22534] = 8'b1111011;
DRAM[22535] = 8'b1111011;
DRAM[22536] = 8'b1111100;
DRAM[22537] = 8'b1111100;
DRAM[22538] = 8'b1111100;
DRAM[22539] = 8'b1111101;
DRAM[22540] = 8'b1111101;
DRAM[22541] = 8'b1111110;
DRAM[22542] = 8'b1111110;
DRAM[22543] = 8'b1111110;
DRAM[22544] = 8'b10000000;
DRAM[22545] = 8'b1111110;
DRAM[22546] = 8'b1111110;
DRAM[22547] = 8'b10000001;
DRAM[22548] = 8'b10000010;
DRAM[22549] = 8'b10000011;
DRAM[22550] = 8'b10001000;
DRAM[22551] = 8'b10001110;
DRAM[22552] = 8'b10011000;
DRAM[22553] = 8'b10100110;
DRAM[22554] = 8'b10111011;
DRAM[22555] = 8'b11010010;
DRAM[22556] = 8'b11100110;
DRAM[22557] = 8'b11110100;
DRAM[22558] = 8'b11111010;
DRAM[22559] = 8'b11111011;
DRAM[22560] = 8'b11101100;
DRAM[22561] = 8'b11101011;
DRAM[22562] = 8'b11100001;
DRAM[22563] = 8'b11101101;
DRAM[22564] = 8'b11111111;
DRAM[22565] = 8'b11100110;
DRAM[22566] = 8'b11010100;
DRAM[22567] = 8'b11101100;
DRAM[22568] = 8'b11100011;
DRAM[22569] = 8'b11101100;
DRAM[22570] = 8'b11010111;
DRAM[22571] = 8'b11010101;
DRAM[22572] = 8'b11101101;
DRAM[22573] = 8'b11011100;
DRAM[22574] = 8'b11001000;
DRAM[22575] = 8'b11100010;
DRAM[22576] = 8'b11010010;
DRAM[22577] = 8'b11001010;
DRAM[22578] = 8'b11101101;
DRAM[22579] = 8'b11010000;
DRAM[22580] = 8'b11101001;
DRAM[22581] = 8'b11101001;
DRAM[22582] = 8'b11000001;
DRAM[22583] = 8'b10110110;
DRAM[22584] = 8'b11011111;
DRAM[22585] = 8'b11011111;
DRAM[22586] = 8'b11110100;
DRAM[22587] = 8'b11001000;
DRAM[22588] = 8'b11001001;
DRAM[22589] = 8'b11101001;
DRAM[22590] = 8'b11001101;
DRAM[22591] = 8'b11011101;
DRAM[22592] = 8'b11110001;
DRAM[22593] = 8'b11100111;
DRAM[22594] = 8'b11100010;
DRAM[22595] = 8'b11101010;
DRAM[22596] = 8'b11110010;
DRAM[22597] = 8'b11101101;
DRAM[22598] = 8'b11011101;
DRAM[22599] = 8'b11010001;
DRAM[22600] = 8'b10111010;
DRAM[22601] = 8'b10011100;
DRAM[22602] = 8'b10101111;
DRAM[22603] = 8'b10011110;
DRAM[22604] = 8'b1110000;
DRAM[22605] = 8'b1011101;
DRAM[22606] = 8'b1011011;
DRAM[22607] = 8'b1110111;
DRAM[22608] = 8'b1110110;
DRAM[22609] = 8'b10000100;
DRAM[22610] = 8'b10001011;
DRAM[22611] = 8'b10010111;
DRAM[22612] = 8'b10110001;
DRAM[22613] = 8'b11000011;
DRAM[22614] = 8'b11000111;
DRAM[22615] = 8'b11001010;
DRAM[22616] = 8'b11101001;
DRAM[22617] = 8'b11011101;
DRAM[22618] = 8'b11010101;
DRAM[22619] = 8'b11011001;
DRAM[22620] = 8'b11011110;
DRAM[22621] = 8'b11011010;
DRAM[22622] = 8'b11010000;
DRAM[22623] = 8'b11001001;
DRAM[22624] = 8'b11001000;
DRAM[22625] = 8'b11001110;
DRAM[22626] = 8'b11010010;
DRAM[22627] = 8'b11001011;
DRAM[22628] = 8'b10111110;
DRAM[22629] = 8'b10110110;
DRAM[22630] = 8'b10111001;
DRAM[22631] = 8'b10111110;
DRAM[22632] = 8'b11001010;
DRAM[22633] = 8'b11000001;
DRAM[22634] = 8'b11001011;
DRAM[22635] = 8'b11001110;
DRAM[22636] = 8'b10111000;
DRAM[22637] = 8'b10110000;
DRAM[22638] = 8'b10111000;
DRAM[22639] = 8'b10110110;
DRAM[22640] = 8'b10111000;
DRAM[22641] = 8'b10111000;
DRAM[22642] = 8'b10111011;
DRAM[22643] = 8'b10111101;
DRAM[22644] = 8'b10110111;
DRAM[22645] = 8'b10110000;
DRAM[22646] = 8'b10110110;
DRAM[22647] = 8'b11000011;
DRAM[22648] = 8'b10110110;
DRAM[22649] = 8'b10100101;
DRAM[22650] = 8'b11000010;
DRAM[22651] = 8'b10111111;
DRAM[22652] = 8'b10110110;
DRAM[22653] = 8'b10101011;
DRAM[22654] = 8'b11000011;
DRAM[22655] = 8'b10110011;
DRAM[22656] = 8'b10101100;
DRAM[22657] = 8'b10101101;
DRAM[22658] = 8'b10111001;
DRAM[22659] = 8'b10100010;
DRAM[22660] = 8'b10111101;
DRAM[22661] = 8'b10101011;
DRAM[22662] = 8'b10111110;
DRAM[22663] = 8'b10100111;
DRAM[22664] = 8'b10101100;
DRAM[22665] = 8'b11000010;
DRAM[22666] = 8'b10100111;
DRAM[22667] = 8'b10111010;
DRAM[22668] = 8'b10100001;
DRAM[22669] = 8'b10111000;
DRAM[22670] = 8'b10101111;
DRAM[22671] = 8'b10101011;
DRAM[22672] = 8'b10100100;
DRAM[22673] = 8'b10100101;
DRAM[22674] = 8'b10110010;
DRAM[22675] = 8'b10101001;
DRAM[22676] = 8'b10100100;
DRAM[22677] = 8'b10100111;
DRAM[22678] = 8'b10011010;
DRAM[22679] = 8'b10011010;
DRAM[22680] = 8'b10011101;
DRAM[22681] = 8'b10100000;
DRAM[22682] = 8'b10110100;
DRAM[22683] = 8'b10110011;
DRAM[22684] = 8'b10011011;
DRAM[22685] = 8'b10110000;
DRAM[22686] = 8'b10100001;
DRAM[22687] = 8'b10101010;
DRAM[22688] = 8'b10111010;
DRAM[22689] = 8'b10010000;
DRAM[22690] = 8'b10001110;
DRAM[22691] = 8'b10100010;
DRAM[22692] = 8'b10100000;
DRAM[22693] = 8'b10101110;
DRAM[22694] = 8'b11000011;
DRAM[22695] = 8'b10111111;
DRAM[22696] = 8'b11001001;
DRAM[22697] = 8'b11001111;
DRAM[22698] = 8'b11010001;
DRAM[22699] = 8'b11001101;
DRAM[22700] = 8'b11001001;
DRAM[22701] = 8'b11000110;
DRAM[22702] = 8'b10111111;
DRAM[22703] = 8'b10110101;
DRAM[22704] = 8'b10111101;
DRAM[22705] = 8'b11001010;
DRAM[22706] = 8'b11001011;
DRAM[22707] = 8'b11001001;
DRAM[22708] = 8'b11010000;
DRAM[22709] = 8'b11010011;
DRAM[22710] = 8'b11010101;
DRAM[22711] = 8'b11011101;
DRAM[22712] = 8'b11100011;
DRAM[22713] = 8'b11011111;
DRAM[22714] = 8'b11011111;
DRAM[22715] = 8'b11010101;
DRAM[22716] = 8'b11000001;
DRAM[22717] = 8'b10110011;
DRAM[22718] = 8'b10100100;
DRAM[22719] = 8'b10001111;
DRAM[22720] = 8'b1101001;
DRAM[22721] = 8'b1011000;
DRAM[22722] = 8'b1010001;
DRAM[22723] = 8'b101111;
DRAM[22724] = 8'b1011111;
DRAM[22725] = 8'b10010101;
DRAM[22726] = 8'b10101110;
DRAM[22727] = 8'b10100010;
DRAM[22728] = 8'b10101011;
DRAM[22729] = 8'b10111000;
DRAM[22730] = 8'b11101110;
DRAM[22731] = 8'b11110100;
DRAM[22732] = 8'b11101011;
DRAM[22733] = 8'b11111100;
DRAM[22734] = 8'b11110100;
DRAM[22735] = 8'b11101011;
DRAM[22736] = 8'b11110010;
DRAM[22737] = 8'b11100110;
DRAM[22738] = 8'b11001001;
DRAM[22739] = 8'b11011011;
DRAM[22740] = 8'b10111101;
DRAM[22741] = 8'b11010001;
DRAM[22742] = 8'b11000000;
DRAM[22743] = 8'b11000001;
DRAM[22744] = 8'b11000111;
DRAM[22745] = 8'b11001010;
DRAM[22746] = 8'b11010000;
DRAM[22747] = 8'b10101010;
DRAM[22748] = 8'b10011110;
DRAM[22749] = 8'b11010101;
DRAM[22750] = 8'b10111010;
DRAM[22751] = 8'b11010011;
DRAM[22752] = 8'b11011000;
DRAM[22753] = 8'b11000000;
DRAM[22754] = 8'b10111101;
DRAM[22755] = 8'b11001100;
DRAM[22756] = 8'b10101101;
DRAM[22757] = 8'b11010001;
DRAM[22758] = 8'b11101001;
DRAM[22759] = 8'b11101010;
DRAM[22760] = 8'b11111110;
DRAM[22761] = 8'b11100111;
DRAM[22762] = 8'b11101101;
DRAM[22763] = 8'b10011100;
DRAM[22764] = 8'b1101100;
DRAM[22765] = 8'b10001000;
DRAM[22766] = 8'b1110000;
DRAM[22767] = 8'b1100100;
DRAM[22768] = 8'b1101010;
DRAM[22769] = 8'b1101010;
DRAM[22770] = 8'b1101010;
DRAM[22771] = 8'b1101001;
DRAM[22772] = 8'b1101001;
DRAM[22773] = 8'b1101000;
DRAM[22774] = 8'b1101000;
DRAM[22775] = 8'b1101000;
DRAM[22776] = 8'b1100111;
DRAM[22777] = 8'b1100111;
DRAM[22778] = 8'b1100110;
DRAM[22779] = 8'b1100101;
DRAM[22780] = 8'b1100100;
DRAM[22781] = 8'b1100100;
DRAM[22782] = 8'b1100011;
DRAM[22783] = 8'b1100011;
DRAM[22784] = 8'b1111001;
DRAM[22785] = 8'b1111001;
DRAM[22786] = 8'b1111010;
DRAM[22787] = 8'b1111010;
DRAM[22788] = 8'b1111010;
DRAM[22789] = 8'b1111011;
DRAM[22790] = 8'b1111011;
DRAM[22791] = 8'b1111011;
DRAM[22792] = 8'b1111100;
DRAM[22793] = 8'b1111100;
DRAM[22794] = 8'b1111101;
DRAM[22795] = 8'b1111101;
DRAM[22796] = 8'b1111101;
DRAM[22797] = 8'b1111110;
DRAM[22798] = 8'b1111110;
DRAM[22799] = 8'b1111110;
DRAM[22800] = 8'b1111111;
DRAM[22801] = 8'b1111110;
DRAM[22802] = 8'b10000000;
DRAM[22803] = 8'b10000011;
DRAM[22804] = 8'b10000010;
DRAM[22805] = 8'b10000000;
DRAM[22806] = 8'b10000011;
DRAM[22807] = 8'b10001010;
DRAM[22808] = 8'b10001110;
DRAM[22809] = 8'b10100010;
DRAM[22810] = 8'b10110100;
DRAM[22811] = 8'b11000100;
DRAM[22812] = 8'b11100010;
DRAM[22813] = 8'b11111101;
DRAM[22814] = 8'b11110111;
DRAM[22815] = 8'b11011110;
DRAM[22816] = 8'b11101101;
DRAM[22817] = 8'b11100010;
DRAM[22818] = 8'b11101010;
DRAM[22819] = 8'b11101010;
DRAM[22820] = 8'b11011101;
DRAM[22821] = 8'b11101011;
DRAM[22822] = 8'b11110000;
DRAM[22823] = 8'b11010010;
DRAM[22824] = 8'b11100000;
DRAM[22825] = 8'b11100110;
DRAM[22826] = 8'b11011000;
DRAM[22827] = 8'b11010011;
DRAM[22828] = 8'b11011101;
DRAM[22829] = 8'b11010000;
DRAM[22830] = 8'b11000011;
DRAM[22831] = 8'b11010100;
DRAM[22832] = 8'b11001010;
DRAM[22833] = 8'b11010101;
DRAM[22834] = 8'b11010000;
DRAM[22835] = 8'b10110110;
DRAM[22836] = 8'b11101010;
DRAM[22837] = 8'b11010110;
DRAM[22838] = 8'b10110011;
DRAM[22839] = 8'b11011111;
DRAM[22840] = 8'b11010011;
DRAM[22841] = 8'b11100010;
DRAM[22842] = 8'b11100111;
DRAM[22843] = 8'b11010100;
DRAM[22844] = 8'b11010011;
DRAM[22845] = 8'b11010100;
DRAM[22846] = 8'b11001111;
DRAM[22847] = 8'b11101011;
DRAM[22848] = 8'b11101001;
DRAM[22849] = 8'b11100100;
DRAM[22850] = 8'b11100110;
DRAM[22851] = 8'b11110001;
DRAM[22852] = 8'b11110110;
DRAM[22853] = 8'b11101011;
DRAM[22854] = 8'b11010110;
DRAM[22855] = 8'b11000111;
DRAM[22856] = 8'b11001000;
DRAM[22857] = 8'b10101100;
DRAM[22858] = 8'b10101111;
DRAM[22859] = 8'b10011010;
DRAM[22860] = 8'b1100111;
DRAM[22861] = 8'b1001101;
DRAM[22862] = 8'b1010110;
DRAM[22863] = 8'b1101101;
DRAM[22864] = 8'b1111011;
DRAM[22865] = 8'b10011100;
DRAM[22866] = 8'b10110010;
DRAM[22867] = 8'b10110110;
DRAM[22868] = 8'b10111001;
DRAM[22869] = 8'b10111101;
DRAM[22870] = 8'b11001010;
DRAM[22871] = 8'b11011101;
DRAM[22872] = 8'b11000110;
DRAM[22873] = 8'b11001110;
DRAM[22874] = 8'b11011010;
DRAM[22875] = 8'b11100000;
DRAM[22876] = 8'b11011001;
DRAM[22877] = 8'b11001110;
DRAM[22878] = 8'b11001011;
DRAM[22879] = 8'b11001110;
DRAM[22880] = 8'b11000111;
DRAM[22881] = 8'b11001100;
DRAM[22882] = 8'b11010000;
DRAM[22883] = 8'b11001101;
DRAM[22884] = 8'b11000110;
DRAM[22885] = 8'b11000001;
DRAM[22886] = 8'b11000011;
DRAM[22887] = 8'b11000111;
DRAM[22888] = 8'b10111111;
DRAM[22889] = 8'b10110101;
DRAM[22890] = 8'b10111000;
DRAM[22891] = 8'b11000001;
DRAM[22892] = 8'b11000001;
DRAM[22893] = 8'b10111101;
DRAM[22894] = 8'b10111001;
DRAM[22895] = 8'b10110001;
DRAM[22896] = 8'b10111001;
DRAM[22897] = 8'b10110000;
DRAM[22898] = 8'b10101111;
DRAM[22899] = 8'b10110101;
DRAM[22900] = 8'b10110100;
DRAM[22901] = 8'b10101101;
DRAM[22902] = 8'b10101110;
DRAM[22903] = 8'b10111000;
DRAM[22904] = 8'b10110110;
DRAM[22905] = 8'b10100010;
DRAM[22906] = 8'b10111010;
DRAM[22907] = 8'b10111100;
DRAM[22908] = 8'b10110101;
DRAM[22909] = 8'b10101001;
DRAM[22910] = 8'b11000001;
DRAM[22911] = 8'b10111001;
DRAM[22912] = 8'b10110010;
DRAM[22913] = 8'b10011101;
DRAM[22914] = 8'b10100110;
DRAM[22915] = 8'b10100001;
DRAM[22916] = 8'b10111111;
DRAM[22917] = 8'b10100100;
DRAM[22918] = 8'b10110100;
DRAM[22919] = 8'b10101110;
DRAM[22920] = 8'b10100000;
DRAM[22921] = 8'b10111000;
DRAM[22922] = 8'b10100010;
DRAM[22923] = 8'b10111000;
DRAM[22924] = 8'b10100001;
DRAM[22925] = 8'b10111000;
DRAM[22926] = 8'b10110011;
DRAM[22927] = 8'b10110001;
DRAM[22928] = 8'b10011000;
DRAM[22929] = 8'b10011010;
DRAM[22930] = 8'b10101000;
DRAM[22931] = 8'b10100010;
DRAM[22932] = 8'b10100000;
DRAM[22933] = 8'b10100110;
DRAM[22934] = 8'b10011011;
DRAM[22935] = 8'b10011110;
DRAM[22936] = 8'b10010001;
DRAM[22937] = 8'b10011100;
DRAM[22938] = 8'b10110010;
DRAM[22939] = 8'b10110010;
DRAM[22940] = 8'b10011011;
DRAM[22941] = 8'b10110000;
DRAM[22942] = 8'b10100010;
DRAM[22943] = 8'b10100111;
DRAM[22944] = 8'b10110111;
DRAM[22945] = 8'b10000010;
DRAM[22946] = 8'b10000101;
DRAM[22947] = 8'b10101100;
DRAM[22948] = 8'b10101110;
DRAM[22949] = 8'b10101000;
DRAM[22950] = 8'b10110101;
DRAM[22951] = 8'b10111100;
DRAM[22952] = 8'b10101110;
DRAM[22953] = 8'b10110011;
DRAM[22954] = 8'b10110110;
DRAM[22955] = 8'b10110111;
DRAM[22956] = 8'b10111110;
DRAM[22957] = 8'b11001000;
DRAM[22958] = 8'b11001101;
DRAM[22959] = 8'b11001101;
DRAM[22960] = 8'b11011011;
DRAM[22961] = 8'b11001111;
DRAM[22962] = 8'b10111010;
DRAM[22963] = 8'b10111101;
DRAM[22964] = 8'b11011011;
DRAM[22965] = 8'b11101011;
DRAM[22966] = 8'b11100000;
DRAM[22967] = 8'b11010101;
DRAM[22968] = 8'b11001111;
DRAM[22969] = 8'b11001000;
DRAM[22970] = 8'b11001010;
DRAM[22971] = 8'b11010000;
DRAM[22972] = 8'b11001111;
DRAM[22973] = 8'b11001011;
DRAM[22974] = 8'b10110110;
DRAM[22975] = 8'b10011000;
DRAM[22976] = 8'b10000010;
DRAM[22977] = 8'b1010110;
DRAM[22978] = 8'b1000010;
DRAM[22979] = 8'b101101;
DRAM[22980] = 8'b1011110;
DRAM[22981] = 8'b10001010;
DRAM[22982] = 8'b10100101;
DRAM[22983] = 8'b10101011;
DRAM[22984] = 8'b10101010;
DRAM[22985] = 8'b10110101;
DRAM[22986] = 8'b11101010;
DRAM[22987] = 8'b11110101;
DRAM[22988] = 8'b11101010;
DRAM[22989] = 8'b11110101;
DRAM[22990] = 8'b11110010;
DRAM[22991] = 8'b11110000;
DRAM[22992] = 8'b11101001;
DRAM[22993] = 8'b11011100;
DRAM[22994] = 8'b11001010;
DRAM[22995] = 8'b11011100;
DRAM[22996] = 8'b11000101;
DRAM[22997] = 8'b11001011;
DRAM[22998] = 8'b10111000;
DRAM[22999] = 8'b10110100;
DRAM[23000] = 8'b11001101;
DRAM[23001] = 8'b11000110;
DRAM[23002] = 8'b11001100;
DRAM[23003] = 8'b11000000;
DRAM[23004] = 8'b10101110;
DRAM[23005] = 8'b11000110;
DRAM[23006] = 8'b10110110;
DRAM[23007] = 8'b11010001;
DRAM[23008] = 8'b11001011;
DRAM[23009] = 8'b11100000;
DRAM[23010] = 8'b10111011;
DRAM[23011] = 8'b10110110;
DRAM[23012] = 8'b10111101;
DRAM[23013] = 8'b11010000;
DRAM[23014] = 8'b11010101;
DRAM[23015] = 8'b11110001;
DRAM[23016] = 8'b11110000;
DRAM[23017] = 8'b11101000;
DRAM[23018] = 8'b11110111;
DRAM[23019] = 8'b10111111;
DRAM[23020] = 8'b10000110;
DRAM[23021] = 8'b10000010;
DRAM[23022] = 8'b1110011;
DRAM[23023] = 8'b1110011;
DRAM[23024] = 8'b1101010;
DRAM[23025] = 8'b1101010;
DRAM[23026] = 8'b1101010;
DRAM[23027] = 8'b1101001;
DRAM[23028] = 8'b1101001;
DRAM[23029] = 8'b1101001;
DRAM[23030] = 8'b1101000;
DRAM[23031] = 8'b1101000;
DRAM[23032] = 8'b1100111;
DRAM[23033] = 8'b1100111;
DRAM[23034] = 8'b1100110;
DRAM[23035] = 8'b1100110;
DRAM[23036] = 8'b1100101;
DRAM[23037] = 8'b1100100;
DRAM[23038] = 8'b1100011;
DRAM[23039] = 8'b1100011;
DRAM[23040] = 8'b1111001;
DRAM[23041] = 8'b1111010;
DRAM[23042] = 8'b1111010;
DRAM[23043] = 8'b1111010;
DRAM[23044] = 8'b1111011;
DRAM[23045] = 8'b1111011;
DRAM[23046] = 8'b1111011;
DRAM[23047] = 8'b1111011;
DRAM[23048] = 8'b1111100;
DRAM[23049] = 8'b1111101;
DRAM[23050] = 8'b1111101;
DRAM[23051] = 8'b1111101;
DRAM[23052] = 8'b1111110;
DRAM[23053] = 8'b1111110;
DRAM[23054] = 8'b1111110;
DRAM[23055] = 8'b1111110;
DRAM[23056] = 8'b1111101;
DRAM[23057] = 8'b1111111;
DRAM[23058] = 8'b10000010;
DRAM[23059] = 8'b10000101;
DRAM[23060] = 8'b10000001;
DRAM[23061] = 8'b1111101;
DRAM[23062] = 8'b10000001;
DRAM[23063] = 8'b10001000;
DRAM[23064] = 8'b10011010;
DRAM[23065] = 8'b10011101;
DRAM[23066] = 8'b10100001;
DRAM[23067] = 8'b10110101;
DRAM[23068] = 8'b11011011;
DRAM[23069] = 8'b11111010;
DRAM[23070] = 8'b11110110;
DRAM[23071] = 8'b11100000;
DRAM[23072] = 8'b11100010;
DRAM[23073] = 8'b11011110;
DRAM[23074] = 8'b11101000;
DRAM[23075] = 8'b11100001;
DRAM[23076] = 8'b11010001;
DRAM[23077] = 8'b11100000;
DRAM[23078] = 8'b11100101;
DRAM[23079] = 8'b11000100;
DRAM[23080] = 8'b11011110;
DRAM[23081] = 8'b11011101;
DRAM[23082] = 8'b11011000;
DRAM[23083] = 8'b11010010;
DRAM[23084] = 8'b11001101;
DRAM[23085] = 8'b11000111;
DRAM[23086] = 8'b11000100;
DRAM[23087] = 8'b11000111;
DRAM[23088] = 8'b11000111;
DRAM[23089] = 8'b11000111;
DRAM[23090] = 8'b11001001;
DRAM[23091] = 8'b11000001;
DRAM[23092] = 8'b11010011;
DRAM[23093] = 8'b11001101;
DRAM[23094] = 8'b11010010;
DRAM[23095] = 8'b11100011;
DRAM[23096] = 8'b10111111;
DRAM[23097] = 8'b11011110;
DRAM[23098] = 8'b11001111;
DRAM[23099] = 8'b11001111;
DRAM[23100] = 8'b11011010;
DRAM[23101] = 8'b11001101;
DRAM[23102] = 8'b11010111;
DRAM[23103] = 8'b11101011;
DRAM[23104] = 8'b11100111;
DRAM[23105] = 8'b11100100;
DRAM[23106] = 8'b11101001;
DRAM[23107] = 8'b11110010;
DRAM[23108] = 8'b11110100;
DRAM[23109] = 8'b11100110;
DRAM[23110] = 8'b11010001;
DRAM[23111] = 8'b11000011;
DRAM[23112] = 8'b10101110;
DRAM[23113] = 8'b10100110;
DRAM[23114] = 8'b10101000;
DRAM[23115] = 8'b10100100;
DRAM[23116] = 8'b1110011;
DRAM[23117] = 8'b1010000;
DRAM[23118] = 8'b1011111;
DRAM[23119] = 8'b1100110;
DRAM[23120] = 8'b1100001;
DRAM[23121] = 8'b1110101;
DRAM[23122] = 8'b10001000;
DRAM[23123] = 8'b10011111;
DRAM[23124] = 8'b10111111;
DRAM[23125] = 8'b11010000;
DRAM[23126] = 8'b11010011;
DRAM[23127] = 8'b11010111;
DRAM[23128] = 8'b11010010;
DRAM[23129] = 8'b11010011;
DRAM[23130] = 8'b11010011;
DRAM[23131] = 8'b11001101;
DRAM[23132] = 8'b11000010;
DRAM[23133] = 8'b10111110;
DRAM[23134] = 8'b11001001;
DRAM[23135] = 8'b11011000;
DRAM[23136] = 8'b11011110;
DRAM[23137] = 8'b11001111;
DRAM[23138] = 8'b11000100;
DRAM[23139] = 8'b11001010;
DRAM[23140] = 8'b11011001;
DRAM[23141] = 8'b11011101;
DRAM[23142] = 8'b11001111;
DRAM[23143] = 8'b10111111;
DRAM[23144] = 8'b11001010;
DRAM[23145] = 8'b11000100;
DRAM[23146] = 8'b10111010;
DRAM[23147] = 8'b10111010;
DRAM[23148] = 8'b11000011;
DRAM[23149] = 8'b11000001;
DRAM[23150] = 8'b10111100;
DRAM[23151] = 8'b10111111;
DRAM[23152] = 8'b11000010;
DRAM[23153] = 8'b10110000;
DRAM[23154] = 8'b10101000;
DRAM[23155] = 8'b10110010;
DRAM[23156] = 8'b10110111;
DRAM[23157] = 8'b10101110;
DRAM[23158] = 8'b10101100;
DRAM[23159] = 8'b10110100;
DRAM[23160] = 8'b10111111;
DRAM[23161] = 8'b10100110;
DRAM[23162] = 8'b10110101;
DRAM[23163] = 8'b10111100;
DRAM[23164] = 8'b10110011;
DRAM[23165] = 8'b10100011;
DRAM[23166] = 8'b10110100;
DRAM[23167] = 8'b10110100;
DRAM[23168] = 8'b10110101;
DRAM[23169] = 8'b10011100;
DRAM[23170] = 8'b10100010;
DRAM[23171] = 8'b10011100;
DRAM[23172] = 8'b10111000;
DRAM[23173] = 8'b10100110;
DRAM[23174] = 8'b10101111;
DRAM[23175] = 8'b10101010;
DRAM[23176] = 8'b10010101;
DRAM[23177] = 8'b10101111;
DRAM[23178] = 8'b10100001;
DRAM[23179] = 8'b10110101;
DRAM[23180] = 8'b10100010;
DRAM[23181] = 8'b10110011;
DRAM[23182] = 8'b10110011;
DRAM[23183] = 8'b10110011;
DRAM[23184] = 8'b10010111;
DRAM[23185] = 8'b10011010;
DRAM[23186] = 8'b10101000;
DRAM[23187] = 8'b10100001;
DRAM[23188] = 8'b10011111;
DRAM[23189] = 8'b10100110;
DRAM[23190] = 8'b10011110;
DRAM[23191] = 8'b10100011;
DRAM[23192] = 8'b10010000;
DRAM[23193] = 8'b10011111;
DRAM[23194] = 8'b10101110;
DRAM[23195] = 8'b10101100;
DRAM[23196] = 8'b10010110;
DRAM[23197] = 8'b10110000;
DRAM[23198] = 8'b10101000;
DRAM[23199] = 8'b10100110;
DRAM[23200] = 8'b10110000;
DRAM[23201] = 8'b10000110;
DRAM[23202] = 8'b10001011;
DRAM[23203] = 8'b10110000;
DRAM[23204] = 8'b10110100;
DRAM[23205] = 8'b10101010;
DRAM[23206] = 8'b10101011;
DRAM[23207] = 8'b10101010;
DRAM[23208] = 8'b10110000;
DRAM[23209] = 8'b10111001;
DRAM[23210] = 8'b11000011;
DRAM[23211] = 8'b11001011;
DRAM[23212] = 8'b11010010;
DRAM[23213] = 8'b11010110;
DRAM[23214] = 8'b11010100;
DRAM[23215] = 8'b11010000;
DRAM[23216] = 8'b11001101;
DRAM[23217] = 8'b11010100;
DRAM[23218] = 8'b11010011;
DRAM[23219] = 8'b11011000;
DRAM[23220] = 8'b11101000;
DRAM[23221] = 8'b11100110;
DRAM[23222] = 8'b11010100;
DRAM[23223] = 8'b11001001;
DRAM[23224] = 8'b11010100;
DRAM[23225] = 8'b11001100;
DRAM[23226] = 8'b11001110;
DRAM[23227] = 8'b11010110;
DRAM[23228] = 8'b11011000;
DRAM[23229] = 8'b11010111;
DRAM[23230] = 8'b11000110;
DRAM[23231] = 8'b10101011;
DRAM[23232] = 8'b10011000;
DRAM[23233] = 8'b1100100;
DRAM[23234] = 8'b1000001;
DRAM[23235] = 8'b101010;
DRAM[23236] = 8'b1010111;
DRAM[23237] = 8'b10001010;
DRAM[23238] = 8'b10100100;
DRAM[23239] = 8'b10101011;
DRAM[23240] = 8'b10101010;
DRAM[23241] = 8'b10110001;
DRAM[23242] = 8'b11100010;
DRAM[23243] = 8'b11110110;
DRAM[23244] = 8'b11101011;
DRAM[23245] = 8'b11101101;
DRAM[23246] = 8'b11101111;
DRAM[23247] = 8'b11110001;
DRAM[23248] = 8'b11101110;
DRAM[23249] = 8'b11011010;
DRAM[23250] = 8'b11010001;
DRAM[23251] = 8'b11011100;
DRAM[23252] = 8'b11010000;
DRAM[23253] = 8'b11001001;
DRAM[23254] = 8'b10111101;
DRAM[23255] = 8'b10110110;
DRAM[23256] = 8'b11000110;
DRAM[23257] = 8'b10110110;
DRAM[23258] = 8'b10111001;
DRAM[23259] = 8'b11001110;
DRAM[23260] = 8'b10111001;
DRAM[23261] = 8'b10101111;
DRAM[23262] = 8'b10101111;
DRAM[23263] = 8'b11000101;
DRAM[23264] = 8'b11000100;
DRAM[23265] = 8'b11101001;
DRAM[23266] = 8'b10111001;
DRAM[23267] = 8'b10101111;
DRAM[23268] = 8'b11000000;
DRAM[23269] = 8'b11000101;
DRAM[23270] = 8'b11001111;
DRAM[23271] = 8'b11101010;
DRAM[23272] = 8'b11101010;
DRAM[23273] = 8'b11100110;
DRAM[23274] = 8'b11100101;
DRAM[23275] = 8'b11001001;
DRAM[23276] = 8'b10010010;
DRAM[23277] = 8'b1101111;
DRAM[23278] = 8'b1101000;
DRAM[23279] = 8'b1101001;
DRAM[23280] = 8'b1101010;
DRAM[23281] = 8'b1101010;
DRAM[23282] = 8'b1101010;
DRAM[23283] = 8'b1101010;
DRAM[23284] = 8'b1101001;
DRAM[23285] = 8'b1101001;
DRAM[23286] = 8'b1101001;
DRAM[23287] = 8'b1101000;
DRAM[23288] = 8'b1101000;
DRAM[23289] = 8'b1101000;
DRAM[23290] = 8'b1100111;
DRAM[23291] = 8'b1100110;
DRAM[23292] = 8'b1100101;
DRAM[23293] = 8'b1100101;
DRAM[23294] = 8'b1100100;
DRAM[23295] = 8'b1100100;
DRAM[23296] = 8'b1111010;
DRAM[23297] = 8'b1111010;
DRAM[23298] = 8'b1111010;
DRAM[23299] = 8'b1111011;
DRAM[23300] = 8'b1111011;
DRAM[23301] = 8'b1111011;
DRAM[23302] = 8'b1111100;
DRAM[23303] = 8'b1111100;
DRAM[23304] = 8'b1111101;
DRAM[23305] = 8'b1111101;
DRAM[23306] = 8'b1111101;
DRAM[23307] = 8'b1111110;
DRAM[23308] = 8'b1111110;
DRAM[23309] = 8'b1111110;
DRAM[23310] = 8'b1111111;
DRAM[23311] = 8'b1111111;
DRAM[23312] = 8'b1111110;
DRAM[23313] = 8'b10000000;
DRAM[23314] = 8'b10000011;
DRAM[23315] = 8'b10000100;
DRAM[23316] = 8'b10000000;
DRAM[23317] = 8'b1111101;
DRAM[23318] = 8'b10000011;
DRAM[23319] = 8'b10001100;
DRAM[23320] = 8'b10100001;
DRAM[23321] = 8'b10010011;
DRAM[23322] = 8'b10011100;
DRAM[23323] = 8'b11000110;
DRAM[23324] = 8'b11101010;
DRAM[23325] = 8'b11110010;
DRAM[23326] = 8'b11101110;
DRAM[23327] = 8'b11101110;
DRAM[23328] = 8'b11001111;
DRAM[23329] = 8'b11011111;
DRAM[23330] = 8'b11011010;
DRAM[23331] = 8'b11011001;
DRAM[23332] = 8'b11011100;
DRAM[23333] = 8'b11000010;
DRAM[23334] = 8'b10110101;
DRAM[23335] = 8'b11001111;
DRAM[23336] = 8'b11100000;
DRAM[23337] = 8'b11010101;
DRAM[23338] = 8'b11010101;
DRAM[23339] = 8'b11010010;
DRAM[23340] = 8'b11000110;
DRAM[23341] = 8'b11001000;
DRAM[23342] = 8'b11001100;
DRAM[23343] = 8'b11000001;
DRAM[23344] = 8'b10111010;
DRAM[23345] = 8'b11000111;
DRAM[23346] = 8'b11010000;
DRAM[23347] = 8'b11001101;
DRAM[23348] = 8'b11001001;
DRAM[23349] = 8'b11010100;
DRAM[23350] = 8'b11100100;
DRAM[23351] = 8'b11001001;
DRAM[23352] = 8'b11000100;
DRAM[23353] = 8'b11011101;
DRAM[23354] = 8'b11000111;
DRAM[23355] = 8'b11000011;
DRAM[23356] = 8'b11011100;
DRAM[23357] = 8'b11010111;
DRAM[23358] = 8'b11010010;
DRAM[23359] = 8'b11011011;
DRAM[23360] = 8'b11101011;
DRAM[23361] = 8'b11100111;
DRAM[23362] = 8'b11101000;
DRAM[23363] = 8'b11101101;
DRAM[23364] = 8'b11101100;
DRAM[23365] = 8'b11011111;
DRAM[23366] = 8'b11001111;
DRAM[23367] = 8'b11000101;
DRAM[23368] = 8'b11010001;
DRAM[23369] = 8'b11000010;
DRAM[23370] = 8'b10100010;
DRAM[23371] = 8'b10001011;
DRAM[23372] = 8'b1010100;
DRAM[23373] = 8'b111001;
DRAM[23374] = 8'b1100101;
DRAM[23375] = 8'b1110001;
DRAM[23376] = 8'b10000110;
DRAM[23377] = 8'b10100000;
DRAM[23378] = 8'b10110010;
DRAM[23379] = 8'b10111000;
DRAM[23380] = 8'b10111010;
DRAM[23381] = 8'b10110101;
DRAM[23382] = 8'b10110111;
DRAM[23383] = 8'b11000011;
DRAM[23384] = 8'b11011000;
DRAM[23385] = 8'b11011000;
DRAM[23386] = 8'b11011111;
DRAM[23387] = 8'b11101000;
DRAM[23388] = 8'b11101000;
DRAM[23389] = 8'b11011100;
DRAM[23390] = 8'b11001101;
DRAM[23391] = 8'b11000100;
DRAM[23392] = 8'b11000000;
DRAM[23393] = 8'b11001111;
DRAM[23394] = 8'b11011010;
DRAM[23395] = 8'b11010001;
DRAM[23396] = 8'b10111110;
DRAM[23397] = 8'b10110100;
DRAM[23398] = 8'b10111100;
DRAM[23399] = 8'b11001010;
DRAM[23400] = 8'b11000001;
DRAM[23401] = 8'b11001111;
DRAM[23402] = 8'b11001011;
DRAM[23403] = 8'b11000110;
DRAM[23404] = 8'b11001011;
DRAM[23405] = 8'b11000010;
DRAM[23406] = 8'b10111011;
DRAM[23407] = 8'b11001001;
DRAM[23408] = 8'b11001100;
DRAM[23409] = 8'b10111000;
DRAM[23410] = 8'b10110000;
DRAM[23411] = 8'b10111001;
DRAM[23412] = 8'b10111101;
DRAM[23413] = 8'b10110101;
DRAM[23414] = 8'b10110100;
DRAM[23415] = 8'b10111100;
DRAM[23416] = 8'b10111110;
DRAM[23417] = 8'b10100110;
DRAM[23418] = 8'b10101110;
DRAM[23419] = 8'b10111101;
DRAM[23420] = 8'b10110100;
DRAM[23421] = 8'b10100011;
DRAM[23422] = 8'b10101001;
DRAM[23423] = 8'b10110000;
DRAM[23424] = 8'b10110000;
DRAM[23425] = 8'b10101011;
DRAM[23426] = 8'b10110100;
DRAM[23427] = 8'b10011010;
DRAM[23428] = 8'b10101100;
DRAM[23429] = 8'b10110001;
DRAM[23430] = 8'b10110001;
DRAM[23431] = 8'b10100000;
DRAM[23432] = 8'b10010101;
DRAM[23433] = 8'b10101101;
DRAM[23434] = 8'b10100101;
DRAM[23435] = 8'b10110101;
DRAM[23436] = 8'b10100100;
DRAM[23437] = 8'b10101100;
DRAM[23438] = 8'b10101110;
DRAM[23439] = 8'b10101101;
DRAM[23440] = 8'b10100000;
DRAM[23441] = 8'b10100010;
DRAM[23442] = 8'b10101110;
DRAM[23443] = 8'b10100011;
DRAM[23444] = 8'b10011110;
DRAM[23445] = 8'b10100011;
DRAM[23446] = 8'b10011011;
DRAM[23447] = 8'b10100000;
DRAM[23448] = 8'b10011010;
DRAM[23449] = 8'b10100101;
DRAM[23450] = 8'b10100110;
DRAM[23451] = 8'b10100011;
DRAM[23452] = 8'b10010100;
DRAM[23453] = 8'b10110001;
DRAM[23454] = 8'b10101110;
DRAM[23455] = 8'b10100011;
DRAM[23456] = 8'b10100101;
DRAM[23457] = 8'b10010110;
DRAM[23458] = 8'b10011010;
DRAM[23459] = 8'b10100110;
DRAM[23460] = 8'b10101001;
DRAM[23461] = 8'b10101100;
DRAM[23462] = 8'b10100011;
DRAM[23463] = 8'b10001101;
DRAM[23464] = 8'b10010100;
DRAM[23465] = 8'b10011110;
DRAM[23466] = 8'b10101111;
DRAM[23467] = 8'b10111111;
DRAM[23468] = 8'b11001100;
DRAM[23469] = 8'b11010100;
DRAM[23470] = 8'b11010110;
DRAM[23471] = 8'b11010101;
DRAM[23472] = 8'b11011011;
DRAM[23473] = 8'b11101000;
DRAM[23474] = 8'b11100100;
DRAM[23475] = 8'b11010100;
DRAM[23476] = 8'b11001101;
DRAM[23477] = 8'b11001100;
DRAM[23478] = 8'b11010010;
DRAM[23479] = 8'b11100001;
DRAM[23480] = 8'b11011000;
DRAM[23481] = 8'b11010100;
DRAM[23482] = 8'b11010110;
DRAM[23483] = 8'b11010010;
DRAM[23484] = 8'b11000111;
DRAM[23485] = 8'b11000110;
DRAM[23486] = 8'b11000100;
DRAM[23487] = 8'b10110111;
DRAM[23488] = 8'b10011000;
DRAM[23489] = 8'b1111010;
DRAM[23490] = 8'b1010110;
DRAM[23491] = 8'b101111;
DRAM[23492] = 8'b1010001;
DRAM[23493] = 8'b10010011;
DRAM[23494] = 8'b10100111;
DRAM[23495] = 8'b10011111;
DRAM[23496] = 8'b10101100;
DRAM[23497] = 8'b10101101;
DRAM[23498] = 8'b11010111;
DRAM[23499] = 8'b11111000;
DRAM[23500] = 8'b11110010;
DRAM[23501] = 8'b11101011;
DRAM[23502] = 8'b11101011;
DRAM[23503] = 8'b11101000;
DRAM[23504] = 8'b11110111;
DRAM[23505] = 8'b11011100;
DRAM[23506] = 8'b11010010;
DRAM[23507] = 8'b11010011;
DRAM[23508] = 8'b11001110;
DRAM[23509] = 8'b11000101;
DRAM[23510] = 8'b11000111;
DRAM[23511] = 8'b11000100;
DRAM[23512] = 8'b10111011;
DRAM[23513] = 8'b10101011;
DRAM[23514] = 8'b10100110;
DRAM[23515] = 8'b11001010;
DRAM[23516] = 8'b10111111;
DRAM[23517] = 8'b10100100;
DRAM[23518] = 8'b10110010;
DRAM[23519] = 8'b10111000;
DRAM[23520] = 8'b11000101;
DRAM[23521] = 8'b11001111;
DRAM[23522] = 8'b10110101;
DRAM[23523] = 8'b10111101;
DRAM[23524] = 8'b10111001;
DRAM[23525] = 8'b10110110;
DRAM[23526] = 8'b11010111;
DRAM[23527] = 8'b11011100;
DRAM[23528] = 8'b11111100;
DRAM[23529] = 8'b11110001;
DRAM[23530] = 8'b11001111;
DRAM[23531] = 8'b10111111;
DRAM[23532] = 8'b10011111;
DRAM[23533] = 8'b1111011;
DRAM[23534] = 8'b1111010;
DRAM[23535] = 8'b1101101;
DRAM[23536] = 8'b1101011;
DRAM[23537] = 8'b1101011;
DRAM[23538] = 8'b1101010;
DRAM[23539] = 8'b1101010;
DRAM[23540] = 8'b1101010;
DRAM[23541] = 8'b1101001;
DRAM[23542] = 8'b1101001;
DRAM[23543] = 8'b1101001;
DRAM[23544] = 8'b1101001;
DRAM[23545] = 8'b1101000;
DRAM[23546] = 8'b1101000;
DRAM[23547] = 8'b1100111;
DRAM[23548] = 8'b1100110;
DRAM[23549] = 8'b1100101;
DRAM[23550] = 8'b1100101;
DRAM[23551] = 8'b1100101;
DRAM[23552] = 8'b1111010;
DRAM[23553] = 8'b1111010;
DRAM[23554] = 8'b1111011;
DRAM[23555] = 8'b1111011;
DRAM[23556] = 8'b1111011;
DRAM[23557] = 8'b1111100;
DRAM[23558] = 8'b1111100;
DRAM[23559] = 8'b1111100;
DRAM[23560] = 8'b1111101;
DRAM[23561] = 8'b1111101;
DRAM[23562] = 8'b1111110;
DRAM[23563] = 8'b1111110;
DRAM[23564] = 8'b1111110;
DRAM[23565] = 8'b1111111;
DRAM[23566] = 8'b1111111;
DRAM[23567] = 8'b1111111;
DRAM[23568] = 8'b10000001;
DRAM[23569] = 8'b10000000;
DRAM[23570] = 8'b10000001;
DRAM[23571] = 8'b10000011;
DRAM[23572] = 8'b10000001;
DRAM[23573] = 8'b10000000;
DRAM[23574] = 8'b10001000;
DRAM[23575] = 8'b10010010;
DRAM[23576] = 8'b10001100;
DRAM[23577] = 8'b10010010;
DRAM[23578] = 8'b10110011;
DRAM[23579] = 8'b11100011;
DRAM[23580] = 8'b11111011;
DRAM[23581] = 8'b11110010;
DRAM[23582] = 8'b11100100;
DRAM[23583] = 8'b11100001;
DRAM[23584] = 8'b11001101;
DRAM[23585] = 8'b11011100;
DRAM[23586] = 8'b11011000;
DRAM[23587] = 8'b11010100;
DRAM[23588] = 8'b11001011;
DRAM[23589] = 8'b10101010;
DRAM[23590] = 8'b10101011;
DRAM[23591] = 8'b11011010;
DRAM[23592] = 8'b11100011;
DRAM[23593] = 8'b11001110;
DRAM[23594] = 8'b11001111;
DRAM[23595] = 8'b11010001;
DRAM[23596] = 8'b11000100;
DRAM[23597] = 8'b11001000;
DRAM[23598] = 8'b11001110;
DRAM[23599] = 8'b10111101;
DRAM[23600] = 8'b10111101;
DRAM[23601] = 8'b11011111;
DRAM[23602] = 8'b11000111;
DRAM[23603] = 8'b11000000;
DRAM[23604] = 8'b11011000;
DRAM[23605] = 8'b11011001;
DRAM[23606] = 8'b11001000;
DRAM[23607] = 8'b11001001;
DRAM[23608] = 8'b11010110;
DRAM[23609] = 8'b11010010;
DRAM[23610] = 8'b11001111;
DRAM[23611] = 8'b11001110;
DRAM[23612] = 8'b11011011;
DRAM[23613] = 8'b11010000;
DRAM[23614] = 8'b10111111;
DRAM[23615] = 8'b11100000;
DRAM[23616] = 8'b11101010;
DRAM[23617] = 8'b11100110;
DRAM[23618] = 8'b11100111;
DRAM[23619] = 8'b11101100;
DRAM[23620] = 8'b11101010;
DRAM[23621] = 8'b11011101;
DRAM[23622] = 8'b11001101;
DRAM[23623] = 8'b11000011;
DRAM[23624] = 8'b10110010;
DRAM[23625] = 8'b10110110;
DRAM[23626] = 8'b10101100;
DRAM[23627] = 8'b10100001;
DRAM[23628] = 8'b1101011;
DRAM[23629] = 8'b1001000;
DRAM[23630] = 8'b1100011;
DRAM[23631] = 8'b1100000;
DRAM[23632] = 8'b1110000;
DRAM[23633] = 8'b10000111;
DRAM[23634] = 8'b10011100;
DRAM[23635] = 8'b10101101;
DRAM[23636] = 8'b10111110;
DRAM[23637] = 8'b11000101;
DRAM[23638] = 8'b11001100;
DRAM[23639] = 8'b11011100;
DRAM[23640] = 8'b11010100;
DRAM[23641] = 8'b11000100;
DRAM[23642] = 8'b10110101;
DRAM[23643] = 8'b10110101;
DRAM[23644] = 8'b10111011;
DRAM[23645] = 8'b11000000;
DRAM[23646] = 8'b11000010;
DRAM[23647] = 8'b11000011;
DRAM[23648] = 8'b10111111;
DRAM[23649] = 8'b10110100;
DRAM[23650] = 8'b10101100;
DRAM[23651] = 8'b10101111;
DRAM[23652] = 8'b10111001;
DRAM[23653] = 8'b10111100;
DRAM[23654] = 8'b10110011;
DRAM[23655] = 8'b10101000;
DRAM[23656] = 8'b10101000;
DRAM[23657] = 8'b11000000;
DRAM[23658] = 8'b11001000;
DRAM[23659] = 8'b11001011;
DRAM[23660] = 8'b11010101;
DRAM[23661] = 8'b11001001;
DRAM[23662] = 8'b10111001;
DRAM[23663] = 8'b10111101;
DRAM[23664] = 8'b11001010;
DRAM[23665] = 8'b10111110;
DRAM[23666] = 8'b10111000;
DRAM[23667] = 8'b10111100;
DRAM[23668] = 8'b10111100;
DRAM[23669] = 8'b10110111;
DRAM[23670] = 8'b10111010;
DRAM[23671] = 8'b11000100;
DRAM[23672] = 8'b10110100;
DRAM[23673] = 8'b10100100;
DRAM[23674] = 8'b10100111;
DRAM[23675] = 8'b10111101;
DRAM[23676] = 8'b10110111;
DRAM[23677] = 8'b10101001;
DRAM[23678] = 8'b10100101;
DRAM[23679] = 8'b10101111;
DRAM[23680] = 8'b10101011;
DRAM[23681] = 8'b10101100;
DRAM[23682] = 8'b10111101;
DRAM[23683] = 8'b10100001;
DRAM[23684] = 8'b10101000;
DRAM[23685] = 8'b10110011;
DRAM[23686] = 8'b10101011;
DRAM[23687] = 8'b10100001;
DRAM[23688] = 8'b10011010;
DRAM[23689] = 8'b10101110;
DRAM[23690] = 8'b10101000;
DRAM[23691] = 8'b10110101;
DRAM[23692] = 8'b10100111;
DRAM[23693] = 8'b10100110;
DRAM[23694] = 8'b10101010;
DRAM[23695] = 8'b10101001;
DRAM[23696] = 8'b10100100;
DRAM[23697] = 8'b10100101;
DRAM[23698] = 8'b10101111;
DRAM[23699] = 8'b10100001;
DRAM[23700] = 8'b10011000;
DRAM[23701] = 8'b10011101;
DRAM[23702] = 8'b10010110;
DRAM[23703] = 8'b10011100;
DRAM[23704] = 8'b10011001;
DRAM[23705] = 8'b10100001;
DRAM[23706] = 8'b10011001;
DRAM[23707] = 8'b10100010;
DRAM[23708] = 8'b10011010;
DRAM[23709] = 8'b10110011;
DRAM[23710] = 8'b10101101;
DRAM[23711] = 8'b10010111;
DRAM[23712] = 8'b10100000;
DRAM[23713] = 8'b10011100;
DRAM[23714] = 8'b10011100;
DRAM[23715] = 8'b10011110;
DRAM[23716] = 8'b10100010;
DRAM[23717] = 8'b10100111;
DRAM[23718] = 8'b10011100;
DRAM[23719] = 8'b10000110;
DRAM[23720] = 8'b10101000;
DRAM[23721] = 8'b10100111;
DRAM[23722] = 8'b10101010;
DRAM[23723] = 8'b10110011;
DRAM[23724] = 8'b11000000;
DRAM[23725] = 8'b11010001;
DRAM[23726] = 8'b11100001;
DRAM[23727] = 8'b11101100;
DRAM[23728] = 8'b11101001;
DRAM[23729] = 8'b11101011;
DRAM[23730] = 8'b11011111;
DRAM[23731] = 8'b11010110;
DRAM[23732] = 8'b11011100;
DRAM[23733] = 8'b11011110;
DRAM[23734] = 8'b11011011;
DRAM[23735] = 8'b11011101;
DRAM[23736] = 8'b11001101;
DRAM[23737] = 8'b11000111;
DRAM[23738] = 8'b11000111;
DRAM[23739] = 8'b11000001;
DRAM[23740] = 8'b10110110;
DRAM[23741] = 8'b10110111;
DRAM[23742] = 8'b10111000;
DRAM[23743] = 8'b10101101;
DRAM[23744] = 8'b10010011;
DRAM[23745] = 8'b10000010;
DRAM[23746] = 8'b1100101;
DRAM[23747] = 8'b1000011;
DRAM[23748] = 8'b1010101;
DRAM[23749] = 8'b10010000;
DRAM[23750] = 8'b10011011;
DRAM[23751] = 8'b10010110;
DRAM[23752] = 8'b10101101;
DRAM[23753] = 8'b10101011;
DRAM[23754] = 8'b11001011;
DRAM[23755] = 8'b11110111;
DRAM[23756] = 8'b11111001;
DRAM[23757] = 8'b11101110;
DRAM[23758] = 8'b11101010;
DRAM[23759] = 8'b11011011;
DRAM[23760] = 8'b11101101;
DRAM[23761] = 8'b11011000;
DRAM[23762] = 8'b11001111;
DRAM[23763] = 8'b11001010;
DRAM[23764] = 8'b11000011;
DRAM[23765] = 8'b10111111;
DRAM[23766] = 8'b11000110;
DRAM[23767] = 8'b11000101;
DRAM[23768] = 8'b10111001;
DRAM[23769] = 8'b10110100;
DRAM[23770] = 8'b10100101;
DRAM[23771] = 8'b10111110;
DRAM[23772] = 8'b11000010;
DRAM[23773] = 8'b10101010;
DRAM[23774] = 8'b10111011;
DRAM[23775] = 8'b10110000;
DRAM[23776] = 8'b10111111;
DRAM[23777] = 8'b10111011;
DRAM[23778] = 8'b10101111;
DRAM[23779] = 8'b10111110;
DRAM[23780] = 8'b11000010;
DRAM[23781] = 8'b10110100;
DRAM[23782] = 8'b11010000;
DRAM[23783] = 8'b11011110;
DRAM[23784] = 8'b11110101;
DRAM[23785] = 8'b11110010;
DRAM[23786] = 8'b10111111;
DRAM[23787] = 8'b10101011;
DRAM[23788] = 8'b10011010;
DRAM[23789] = 8'b10000010;
DRAM[23790] = 8'b10000111;
DRAM[23791] = 8'b1110001;
DRAM[23792] = 8'b1101011;
DRAM[23793] = 8'b1101011;
DRAM[23794] = 8'b1101011;
DRAM[23795] = 8'b1101010;
DRAM[23796] = 8'b1101010;
DRAM[23797] = 8'b1101010;
DRAM[23798] = 8'b1101001;
DRAM[23799] = 8'b1101001;
DRAM[23800] = 8'b1101001;
DRAM[23801] = 8'b1101001;
DRAM[23802] = 8'b1101001;
DRAM[23803] = 8'b1101000;
DRAM[23804] = 8'b1100111;
DRAM[23805] = 8'b1100110;
DRAM[23806] = 8'b1100110;
DRAM[23807] = 8'b1100101;
DRAM[23808] = 8'b1111011;
DRAM[23809] = 8'b1111011;
DRAM[23810] = 8'b1111011;
DRAM[23811] = 8'b1111011;
DRAM[23812] = 8'b1111100;
DRAM[23813] = 8'b1111100;
DRAM[23814] = 8'b1111100;
DRAM[23815] = 8'b1111101;
DRAM[23816] = 8'b1111110;
DRAM[23817] = 8'b1111110;
DRAM[23818] = 8'b1111110;
DRAM[23819] = 8'b1111110;
DRAM[23820] = 8'b1111111;
DRAM[23821] = 8'b1111111;
DRAM[23822] = 8'b1111111;
DRAM[23823] = 8'b10000000;
DRAM[23824] = 8'b10000010;
DRAM[23825] = 8'b1111111;
DRAM[23826] = 8'b10000000;
DRAM[23827] = 8'b10000011;
DRAM[23828] = 8'b10000100;
DRAM[23829] = 8'b10000100;
DRAM[23830] = 8'b10001010;
DRAM[23831] = 8'b10010001;
DRAM[23832] = 8'b10000011;
DRAM[23833] = 8'b10100001;
DRAM[23834] = 8'b11000010;
DRAM[23835] = 8'b11010110;
DRAM[23836] = 8'b11100110;
DRAM[23837] = 8'b11101111;
DRAM[23838] = 8'b11100111;
DRAM[23839] = 8'b11010110;
DRAM[23840] = 8'b11011000;
DRAM[23841] = 8'b11010101;
DRAM[23842] = 8'b11011110;
DRAM[23843] = 8'b11001011;
DRAM[23844] = 8'b10100011;
DRAM[23845] = 8'b10101100;
DRAM[23846] = 8'b11010000;
DRAM[23847] = 8'b11010110;
DRAM[23848] = 8'b11011101;
DRAM[23849] = 8'b11000110;
DRAM[23850] = 8'b11000110;
DRAM[23851] = 8'b11001101;
DRAM[23852] = 8'b11000011;
DRAM[23853] = 8'b11000010;
DRAM[23854] = 8'b11001000;
DRAM[23855] = 8'b11000000;
DRAM[23856] = 8'b11100110;
DRAM[23857] = 8'b11010001;
DRAM[23858] = 8'b11000000;
DRAM[23859] = 8'b11010001;
DRAM[23860] = 8'b11010100;
DRAM[23861] = 8'b11010010;
DRAM[23862] = 8'b11000100;
DRAM[23863] = 8'b11010100;
DRAM[23864] = 8'b11001011;
DRAM[23865] = 8'b10110110;
DRAM[23866] = 8'b11001100;
DRAM[23867] = 8'b11100000;
DRAM[23868] = 8'b11010101;
DRAM[23869] = 8'b10110111;
DRAM[23870] = 8'b10111100;
DRAM[23871] = 8'b11111101;
DRAM[23872] = 8'b11100010;
DRAM[23873] = 8'b11100000;
DRAM[23874] = 8'b11100100;
DRAM[23875] = 8'b11101101;
DRAM[23876] = 8'b11101110;
DRAM[23877] = 8'b11011111;
DRAM[23878] = 8'b11001010;
DRAM[23879] = 8'b10111011;
DRAM[23880] = 8'b10101011;
DRAM[23881] = 8'b10101001;
DRAM[23882] = 8'b10100010;
DRAM[23883] = 8'b10001101;
DRAM[23884] = 8'b1011110;
DRAM[23885] = 8'b1010010;
DRAM[23886] = 8'b1110101;
DRAM[23887] = 8'b10000000;
DRAM[23888] = 8'b10001001;
DRAM[23889] = 8'b10001011;
DRAM[23890] = 8'b10001110;
DRAM[23891] = 8'b10100010;
DRAM[23892] = 8'b11000000;
DRAM[23893] = 8'b11001000;
DRAM[23894] = 8'b11000000;
DRAM[23895] = 8'b11000000;
DRAM[23896] = 8'b11001100;
DRAM[23897] = 8'b11001111;
DRAM[23898] = 8'b11010111;
DRAM[23899] = 8'b11011101;
DRAM[23900] = 8'b11011001;
DRAM[23901] = 8'b11001101;
DRAM[23902] = 8'b11000100;
DRAM[23903] = 8'b11000001;
DRAM[23904] = 8'b10110011;
DRAM[23905] = 8'b10110110;
DRAM[23906] = 8'b10111000;
DRAM[23907] = 8'b10111000;
DRAM[23908] = 8'b10111000;
DRAM[23909] = 8'b10111010;
DRAM[23910] = 8'b10111111;
DRAM[23911] = 8'b11000100;
DRAM[23912] = 8'b11000001;
DRAM[23913] = 8'b11000010;
DRAM[23914] = 8'b10111010;
DRAM[23915] = 8'b10111010;
DRAM[23916] = 8'b11000111;
DRAM[23917] = 8'b11001001;
DRAM[23918] = 8'b10111101;
DRAM[23919] = 8'b10110101;
DRAM[23920] = 8'b10111101;
DRAM[23921] = 8'b10111011;
DRAM[23922] = 8'b10110111;
DRAM[23923] = 8'b10110011;
DRAM[23924] = 8'b10110000;
DRAM[23925] = 8'b10110011;
DRAM[23926] = 8'b10111010;
DRAM[23927] = 8'b11000010;
DRAM[23928] = 8'b10111010;
DRAM[23929] = 8'b10110001;
DRAM[23930] = 8'b10101010;
DRAM[23931] = 8'b10111101;
DRAM[23932] = 8'b10110100;
DRAM[23933] = 8'b10101000;
DRAM[23934] = 8'b10011000;
DRAM[23935] = 8'b10011111;
DRAM[23936] = 8'b10101010;
DRAM[23937] = 8'b10011110;
DRAM[23938] = 8'b10110100;
DRAM[23939] = 8'b10101000;
DRAM[23940] = 8'b10101000;
DRAM[23941] = 8'b10101011;
DRAM[23942] = 8'b10011100;
DRAM[23943] = 8'b10101010;
DRAM[23944] = 8'b10011110;
DRAM[23945] = 8'b10101101;
DRAM[23946] = 8'b10101000;
DRAM[23947] = 8'b10110010;
DRAM[23948] = 8'b10101010;
DRAM[23949] = 8'b10100100;
DRAM[23950] = 8'b10101010;
DRAM[23951] = 8'b10100110;
DRAM[23952] = 8'b10100110;
DRAM[23953] = 8'b10100110;
DRAM[23954] = 8'b10110000;
DRAM[23955] = 8'b10100010;
DRAM[23956] = 8'b10011010;
DRAM[23957] = 8'b10011111;
DRAM[23958] = 8'b10011011;
DRAM[23959] = 8'b10100101;
DRAM[23960] = 8'b10001110;
DRAM[23961] = 8'b10010110;
DRAM[23962] = 8'b10001111;
DRAM[23963] = 8'b10100111;
DRAM[23964] = 8'b10100011;
DRAM[23965] = 8'b10101111;
DRAM[23966] = 8'b10100100;
DRAM[23967] = 8'b10001000;
DRAM[23968] = 8'b10100001;
DRAM[23969] = 8'b10011000;
DRAM[23970] = 8'b10010110;
DRAM[23971] = 8'b10100001;
DRAM[23972] = 8'b10101000;
DRAM[23973] = 8'b10100010;
DRAM[23974] = 8'b10011011;
DRAM[23975] = 8'b10011011;
DRAM[23976] = 8'b10011101;
DRAM[23977] = 8'b10011001;
DRAM[23978] = 8'b10011000;
DRAM[23979] = 8'b10011110;
DRAM[23980] = 8'b10100111;
DRAM[23981] = 8'b10110010;
DRAM[23982] = 8'b11000000;
DRAM[23983] = 8'b11001100;
DRAM[23984] = 8'b11010011;
DRAM[23985] = 8'b11100000;
DRAM[23986] = 8'b11100111;
DRAM[23987] = 8'b11101110;
DRAM[23988] = 8'b11111011;
DRAM[23989] = 8'b11110110;
DRAM[23990] = 8'b11100010;
DRAM[23991] = 8'b11010111;
DRAM[23992] = 8'b11011011;
DRAM[23993] = 8'b11001100;
DRAM[23994] = 8'b11000101;
DRAM[23995] = 8'b11000011;
DRAM[23996] = 8'b11000001;
DRAM[23997] = 8'b11000010;
DRAM[23998] = 8'b10110110;
DRAM[23999] = 8'b10011110;
DRAM[24000] = 8'b10010100;
DRAM[24001] = 8'b1111110;
DRAM[24002] = 8'b1100110;
DRAM[24003] = 8'b1011001;
DRAM[24004] = 8'b1011100;
DRAM[24005] = 8'b10000011;
DRAM[24006] = 8'b10001000;
DRAM[24007] = 8'b10011000;
DRAM[24008] = 8'b10101011;
DRAM[24009] = 8'b10101010;
DRAM[24010] = 8'b11000010;
DRAM[24011] = 8'b11110011;
DRAM[24012] = 8'b11111100;
DRAM[24013] = 8'b11110010;
DRAM[24014] = 8'b11101111;
DRAM[24015] = 8'b11010101;
DRAM[24016] = 8'b11011101;
DRAM[24017] = 8'b11011001;
DRAM[24018] = 8'b11010100;
DRAM[24019] = 8'b11010001;
DRAM[24020] = 8'b10111110;
DRAM[24021] = 8'b11000011;
DRAM[24022] = 8'b11000011;
DRAM[24023] = 8'b10111111;
DRAM[24024] = 8'b10110110;
DRAM[24025] = 8'b11000000;
DRAM[24026] = 8'b10101101;
DRAM[24027] = 8'b10101100;
DRAM[24028] = 8'b10111111;
DRAM[24029] = 8'b10101101;
DRAM[24030] = 8'b10110110;
DRAM[24031] = 8'b10101010;
DRAM[24032] = 8'b10110001;
DRAM[24033] = 8'b10111001;
DRAM[24034] = 8'b10101101;
DRAM[24035] = 8'b10101000;
DRAM[24036] = 8'b11010001;
DRAM[24037] = 8'b11000000;
DRAM[24038] = 8'b10111110;
DRAM[24039] = 8'b11101001;
DRAM[24040] = 8'b11100110;
DRAM[24041] = 8'b11110010;
DRAM[24042] = 8'b11000101;
DRAM[24043] = 8'b10100010;
DRAM[24044] = 8'b10001010;
DRAM[24045] = 8'b1110011;
DRAM[24046] = 8'b1110101;
DRAM[24047] = 8'b1100110;
DRAM[24048] = 8'b1101100;
DRAM[24049] = 8'b1101011;
DRAM[24050] = 8'b1101011;
DRAM[24051] = 8'b1101011;
DRAM[24052] = 8'b1101010;
DRAM[24053] = 8'b1101010;
DRAM[24054] = 8'b1101010;
DRAM[24055] = 8'b1101010;
DRAM[24056] = 8'b1101010;
DRAM[24057] = 8'b1101010;
DRAM[24058] = 8'b1101001;
DRAM[24059] = 8'b1101001;
DRAM[24060] = 8'b1101000;
DRAM[24061] = 8'b1100111;
DRAM[24062] = 8'b1100110;
DRAM[24063] = 8'b1100110;
DRAM[24064] = 8'b1111011;
DRAM[24065] = 8'b1111011;
DRAM[24066] = 8'b1111011;
DRAM[24067] = 8'b1111100;
DRAM[24068] = 8'b1111100;
DRAM[24069] = 8'b1111100;
DRAM[24070] = 8'b1111101;
DRAM[24071] = 8'b1111101;
DRAM[24072] = 8'b1111110;
DRAM[24073] = 8'b1111110;
DRAM[24074] = 8'b1111110;
DRAM[24075] = 8'b1111111;
DRAM[24076] = 8'b1111111;
DRAM[24077] = 8'b1111111;
DRAM[24078] = 8'b10000000;
DRAM[24079] = 8'b10000000;
DRAM[24080] = 8'b10000010;
DRAM[24081] = 8'b1111110;
DRAM[24082] = 8'b1111111;
DRAM[24083] = 8'b10000100;
DRAM[24084] = 8'b10001000;
DRAM[24085] = 8'b10000111;
DRAM[24086] = 8'b10000111;
DRAM[24087] = 8'b10001000;
DRAM[24088] = 8'b10001100;
DRAM[24089] = 8'b10100011;
DRAM[24090] = 8'b10110011;
DRAM[24091] = 8'b10111010;
DRAM[24092] = 8'b11001101;
DRAM[24093] = 8'b11100111;
DRAM[24094] = 8'b11101011;
DRAM[24095] = 8'b11011101;
DRAM[24096] = 8'b11010111;
DRAM[24097] = 8'b11010110;
DRAM[24098] = 8'b11010101;
DRAM[24099] = 8'b10110111;
DRAM[24100] = 8'b10011110;
DRAM[24101] = 8'b11000001;
DRAM[24102] = 8'b11100010;
DRAM[24103] = 8'b11010001;
DRAM[24104] = 8'b11001011;
DRAM[24105] = 8'b10111010;
DRAM[24106] = 8'b10111110;
DRAM[24107] = 8'b11001010;
DRAM[24108] = 8'b11000011;
DRAM[24109] = 8'b10111011;
DRAM[24110] = 8'b11000101;
DRAM[24111] = 8'b11010001;
DRAM[24112] = 8'b11101110;
DRAM[24113] = 8'b10110010;
DRAM[24114] = 8'b11000100;
DRAM[24115] = 8'b11100110;
DRAM[24116] = 8'b11001001;
DRAM[24117] = 8'b11010100;
DRAM[24118] = 8'b11000111;
DRAM[24119] = 8'b11001011;
DRAM[24120] = 8'b10111100;
DRAM[24121] = 8'b10111000;
DRAM[24122] = 8'b11001011;
DRAM[24123] = 8'b11100111;
DRAM[24124] = 8'b11001011;
DRAM[24125] = 8'b10101110;
DRAM[24126] = 8'b11010111;
DRAM[24127] = 8'b11111111;
DRAM[24128] = 8'b11011111;
DRAM[24129] = 8'b11011010;
DRAM[24130] = 8'b11011100;
DRAM[24131] = 8'b11100110;
DRAM[24132] = 8'b11101010;
DRAM[24133] = 8'b11011110;
DRAM[24134] = 8'b11001000;
DRAM[24135] = 8'b10111001;
DRAM[24136] = 8'b10101011;
DRAM[24137] = 8'b10101001;
DRAM[24138] = 8'b10110111;
DRAM[24139] = 8'b10011001;
DRAM[24140] = 8'b1100011;
DRAM[24141] = 8'b1010101;
DRAM[24142] = 8'b1011100;
DRAM[24143] = 8'b1100100;
DRAM[24144] = 8'b10001101;
DRAM[24145] = 8'b10100101;
DRAM[24146] = 8'b10111001;
DRAM[24147] = 8'b11000011;
DRAM[24148] = 8'b11000100;
DRAM[24149] = 8'b10111101;
DRAM[24150] = 8'b11000101;
DRAM[24151] = 8'b11011100;
DRAM[24152] = 8'b11011100;
DRAM[24153] = 8'b11011000;
DRAM[24154] = 8'b11010100;
DRAM[24155] = 8'b11001110;
DRAM[24156] = 8'b11000110;
DRAM[24157] = 8'b11000001;
DRAM[24158] = 8'b11000110;
DRAM[24159] = 8'b11001111;
DRAM[24160] = 8'b11010110;
DRAM[24161] = 8'b11000111;
DRAM[24162] = 8'b10111010;
DRAM[24163] = 8'b10111111;
DRAM[24164] = 8'b11001111;
DRAM[24165] = 8'b11011000;
DRAM[24166] = 8'b11010011;
DRAM[24167] = 8'b11001001;
DRAM[24168] = 8'b11100000;
DRAM[24169] = 8'b11001111;
DRAM[24170] = 8'b11000001;
DRAM[24171] = 8'b10111001;
DRAM[24172] = 8'b10111001;
DRAM[24173] = 8'b11000100;
DRAM[24174] = 8'b11000110;
DRAM[24175] = 8'b10111010;
DRAM[24176] = 8'b10110001;
DRAM[24177] = 8'b10110110;
DRAM[24178] = 8'b10110010;
DRAM[24179] = 8'b10100111;
DRAM[24180] = 8'b10100111;
DRAM[24181] = 8'b10110011;
DRAM[24182] = 8'b10111100;
DRAM[24183] = 8'b10111011;
DRAM[24184] = 8'b11000010;
DRAM[24185] = 8'b10111110;
DRAM[24186] = 8'b10101110;
DRAM[24187] = 8'b10111001;
DRAM[24188] = 8'b10101110;
DRAM[24189] = 8'b10101000;
DRAM[24190] = 8'b10010000;
DRAM[24191] = 8'b10010100;
DRAM[24192] = 8'b10101011;
DRAM[24193] = 8'b10011011;
DRAM[24194] = 8'b10101110;
DRAM[24195] = 8'b10100010;
DRAM[24196] = 8'b10100000;
DRAM[24197] = 8'b10101100;
DRAM[24198] = 8'b10010110;
DRAM[24199] = 8'b10100101;
DRAM[24200] = 8'b10100101;
DRAM[24201] = 8'b10101101;
DRAM[24202] = 8'b10101000;
DRAM[24203] = 8'b10101110;
DRAM[24204] = 8'b10101011;
DRAM[24205] = 8'b10100000;
DRAM[24206] = 8'b10100111;
DRAM[24207] = 8'b10100001;
DRAM[24208] = 8'b10100100;
DRAM[24209] = 8'b10100110;
DRAM[24210] = 8'b10110001;
DRAM[24211] = 8'b10100011;
DRAM[24212] = 8'b10011100;
DRAM[24213] = 8'b10100100;
DRAM[24214] = 8'b10100011;
DRAM[24215] = 8'b10101110;
DRAM[24216] = 8'b10010010;
DRAM[24217] = 8'b10011000;
DRAM[24218] = 8'b10001110;
DRAM[24219] = 8'b10101100;
DRAM[24220] = 8'b10100001;
DRAM[24221] = 8'b10100000;
DRAM[24222] = 8'b10011010;
DRAM[24223] = 8'b10000100;
DRAM[24224] = 8'b10010001;
DRAM[24225] = 8'b10010010;
DRAM[24226] = 8'b10010000;
DRAM[24227] = 8'b10010110;
DRAM[24228] = 8'b10011111;
DRAM[24229] = 8'b10011110;
DRAM[24230] = 8'b10011100;
DRAM[24231] = 8'b10100010;
DRAM[24232] = 8'b10001001;
DRAM[24233] = 8'b10001000;
DRAM[24234] = 8'b10001110;
DRAM[24235] = 8'b10011100;
DRAM[24236] = 8'b10101001;
DRAM[24237] = 8'b10110010;
DRAM[24238] = 8'b10111110;
DRAM[24239] = 8'b11001001;
DRAM[24240] = 8'b11001110;
DRAM[24241] = 8'b11011111;
DRAM[24242] = 8'b11100100;
DRAM[24243] = 8'b11100010;
DRAM[24244] = 8'b11100111;
DRAM[24245] = 8'b11101001;
DRAM[24246] = 8'b11101011;
DRAM[24247] = 8'b11110100;
DRAM[24248] = 8'b11110010;
DRAM[24249] = 8'b11100001;
DRAM[24250] = 8'b11010110;
DRAM[24251] = 8'b11010001;
DRAM[24252] = 8'b11001100;
DRAM[24253] = 8'b11001101;
DRAM[24254] = 8'b11000001;
DRAM[24255] = 8'b10101001;
DRAM[24256] = 8'b10011001;
DRAM[24257] = 8'b10000011;
DRAM[24258] = 8'b1100111;
DRAM[24259] = 8'b1011010;
DRAM[24260] = 8'b1010111;
DRAM[24261] = 8'b10000001;
DRAM[24262] = 8'b10000110;
DRAM[24263] = 8'b10011001;
DRAM[24264] = 8'b10100101;
DRAM[24265] = 8'b10101010;
DRAM[24266] = 8'b10111110;
DRAM[24267] = 8'b11101101;
DRAM[24268] = 8'b11111000;
DRAM[24269] = 8'b11110100;
DRAM[24270] = 8'b11111001;
DRAM[24271] = 8'b11011010;
DRAM[24272] = 8'b11010111;
DRAM[24273] = 8'b11100101;
DRAM[24274] = 8'b11011110;
DRAM[24275] = 8'b11011011;
DRAM[24276] = 8'b10111000;
DRAM[24277] = 8'b11001010;
DRAM[24278] = 8'b11000011;
DRAM[24279] = 8'b10111100;
DRAM[24280] = 8'b10101010;
DRAM[24281] = 8'b10111111;
DRAM[24282] = 8'b10110001;
DRAM[24283] = 8'b10011101;
DRAM[24284] = 8'b10111011;
DRAM[24285] = 8'b10101001;
DRAM[24286] = 8'b10100111;
DRAM[24287] = 8'b10101101;
DRAM[24288] = 8'b10101100;
DRAM[24289] = 8'b10101000;
DRAM[24290] = 8'b10110010;
DRAM[24291] = 8'b10010111;
DRAM[24292] = 8'b10111111;
DRAM[24293] = 8'b11001011;
DRAM[24294] = 8'b11000010;
DRAM[24295] = 8'b11100001;
DRAM[24296] = 8'b11101111;
DRAM[24297] = 8'b11111000;
DRAM[24298] = 8'b11010011;
DRAM[24299] = 8'b10101000;
DRAM[24300] = 8'b10001101;
DRAM[24301] = 8'b1110101;
DRAM[24302] = 8'b1101101;
DRAM[24303] = 8'b1101110;
DRAM[24304] = 8'b1101100;
DRAM[24305] = 8'b1101100;
DRAM[24306] = 8'b1101011;
DRAM[24307] = 8'b1101011;
DRAM[24308] = 8'b1101011;
DRAM[24309] = 8'b1101010;
DRAM[24310] = 8'b1101010;
DRAM[24311] = 8'b1101010;
DRAM[24312] = 8'b1101011;
DRAM[24313] = 8'b1101011;
DRAM[24314] = 8'b1101010;
DRAM[24315] = 8'b1101001;
DRAM[24316] = 8'b1101000;
DRAM[24317] = 8'b1101000;
DRAM[24318] = 8'b1100111;
DRAM[24319] = 8'b1100111;
DRAM[24320] = 8'b1111011;
DRAM[24321] = 8'b1111011;
DRAM[24322] = 8'b1111011;
DRAM[24323] = 8'b1111100;
DRAM[24324] = 8'b1111100;
DRAM[24325] = 8'b1111101;
DRAM[24326] = 8'b1111101;
DRAM[24327] = 8'b1111101;
DRAM[24328] = 8'b1111110;
DRAM[24329] = 8'b1111110;
DRAM[24330] = 8'b1111110;
DRAM[24331] = 8'b1111111;
DRAM[24332] = 8'b1111111;
DRAM[24333] = 8'b10000000;
DRAM[24334] = 8'b10000000;
DRAM[24335] = 8'b10000000;
DRAM[24336] = 8'b10000001;
DRAM[24337] = 8'b1111101;
DRAM[24338] = 8'b1111110;
DRAM[24339] = 8'b10000110;
DRAM[24340] = 8'b10001100;
DRAM[24341] = 8'b10001000;
DRAM[24342] = 8'b10000010;
DRAM[24343] = 8'b1111111;
DRAM[24344] = 8'b10001110;
DRAM[24345] = 8'b10010010;
DRAM[24346] = 8'b10011111;
DRAM[24347] = 8'b10110111;
DRAM[24348] = 8'b11010011;
DRAM[24349] = 8'b11100101;
DRAM[24350] = 8'b11100110;
DRAM[24351] = 8'b11100000;
DRAM[24352] = 8'b11001011;
DRAM[24353] = 8'b11011101;
DRAM[24354] = 8'b11000001;
DRAM[24355] = 8'b10100100;
DRAM[24356] = 8'b10111011;
DRAM[24357] = 8'b11010011;
DRAM[24358] = 8'b11010010;
DRAM[24359] = 8'b11010011;
DRAM[24360] = 8'b10111010;
DRAM[24361] = 8'b10110000;
DRAM[24362] = 8'b10111000;
DRAM[24363] = 8'b11001001;
DRAM[24364] = 8'b11000101;
DRAM[24365] = 8'b10111001;
DRAM[24366] = 8'b11001000;
DRAM[24367] = 8'b11100101;
DRAM[24368] = 8'b11000000;
DRAM[24369] = 8'b10110100;
DRAM[24370] = 8'b11000110;
DRAM[24371] = 8'b11010111;
DRAM[24372] = 8'b11010111;
DRAM[24373] = 8'b11100000;
DRAM[24374] = 8'b10101000;
DRAM[24375] = 8'b10111101;
DRAM[24376] = 8'b11000110;
DRAM[24377] = 8'b11011110;
DRAM[24378] = 8'b11011000;
DRAM[24379] = 8'b11101000;
DRAM[24380] = 8'b11000101;
DRAM[24381] = 8'b10110111;
DRAM[24382] = 8'b11110011;
DRAM[24383] = 8'b11100010;
DRAM[24384] = 8'b11100011;
DRAM[24385] = 8'b11011000;
DRAM[24386] = 8'b11010011;
DRAM[24387] = 8'b11011010;
DRAM[24388] = 8'b11100001;
DRAM[24389] = 8'b11011010;
DRAM[24390] = 8'b11001010;
DRAM[24391] = 8'b10111101;
DRAM[24392] = 8'b10110111;
DRAM[24393] = 8'b10100111;
DRAM[24394] = 8'b10110001;
DRAM[24395] = 8'b10000011;
DRAM[24396] = 8'b1001111;
DRAM[24397] = 8'b1010100;
DRAM[24398] = 8'b1100010;
DRAM[24399] = 8'b1111001;
DRAM[24400] = 8'b1111001;
DRAM[24401] = 8'b10000111;
DRAM[24402] = 8'b10010101;
DRAM[24403] = 8'b10100110;
DRAM[24404] = 8'b10110100;
DRAM[24405] = 8'b10110001;
DRAM[24406] = 8'b10110000;
DRAM[24407] = 8'b10111100;
DRAM[24408] = 8'b11001011;
DRAM[24409] = 8'b11001000;
DRAM[24410] = 8'b11001000;
DRAM[24411] = 8'b11001101;
DRAM[24412] = 8'b11001110;
DRAM[24413] = 8'b11001010;
DRAM[24414] = 8'b11000111;
DRAM[24415] = 8'b11000111;
DRAM[24416] = 8'b11010011;
DRAM[24417] = 8'b11010110;
DRAM[24418] = 8'b11010110;
DRAM[24419] = 8'b11001101;
DRAM[24420] = 8'b11000010;
DRAM[24421] = 8'b11000000;
DRAM[24422] = 8'b11001001;
DRAM[24423] = 8'b11010011;
DRAM[24424] = 8'b11001111;
DRAM[24425] = 8'b11001010;
DRAM[24426] = 8'b11010010;
DRAM[24427] = 8'b11010000;
DRAM[24428] = 8'b11000001;
DRAM[24429] = 8'b11000110;
DRAM[24430] = 8'b11001100;
DRAM[24431] = 8'b10111101;
DRAM[24432] = 8'b10101101;
DRAM[24433] = 8'b10110101;
DRAM[24434] = 8'b10110000;
DRAM[24435] = 8'b10100001;
DRAM[24436] = 8'b10100100;
DRAM[24437] = 8'b10110111;
DRAM[24438] = 8'b11000000;
DRAM[24439] = 8'b10111000;
DRAM[24440] = 8'b10111010;
DRAM[24441] = 8'b10111100;
DRAM[24442] = 8'b10101000;
DRAM[24443] = 8'b10110011;
DRAM[24444] = 8'b10101011;
DRAM[24445] = 8'b10101111;
DRAM[24446] = 8'b10011000;
DRAM[24447] = 8'b10011101;
DRAM[24448] = 8'b10101010;
DRAM[24449] = 8'b10100110;
DRAM[24450] = 8'b10110011;
DRAM[24451] = 8'b10010100;
DRAM[24452] = 8'b10010010;
DRAM[24453] = 8'b10110100;
DRAM[24454] = 8'b10011001;
DRAM[24455] = 8'b10010110;
DRAM[24456] = 8'b10101011;
DRAM[24457] = 8'b10101111;
DRAM[24458] = 8'b10101000;
DRAM[24459] = 8'b10101011;
DRAM[24460] = 8'b10101010;
DRAM[24461] = 8'b10011100;
DRAM[24462] = 8'b10100010;
DRAM[24463] = 8'b10011010;
DRAM[24464] = 8'b10011111;
DRAM[24465] = 8'b10100001;
DRAM[24466] = 8'b10101100;
DRAM[24467] = 8'b10011110;
DRAM[24468] = 8'b10010111;
DRAM[24469] = 8'b10100000;
DRAM[24470] = 8'b10100001;
DRAM[24471] = 8'b10101101;
DRAM[24472] = 8'b10100001;
DRAM[24473] = 8'b10100100;
DRAM[24474] = 8'b10010010;
DRAM[24475] = 8'b10101011;
DRAM[24476] = 8'b10011000;
DRAM[24477] = 8'b10010000;
DRAM[24478] = 8'b10010011;
DRAM[24479] = 8'b10001000;
DRAM[24480] = 8'b1110100;
DRAM[24481] = 8'b10001100;
DRAM[24482] = 8'b10001100;
DRAM[24483] = 8'b1111101;
DRAM[24484] = 8'b10000111;
DRAM[24485] = 8'b10011000;
DRAM[24486] = 8'b10010111;
DRAM[24487] = 8'b10001111;
DRAM[24488] = 8'b10001111;
DRAM[24489] = 8'b10000101;
DRAM[24490] = 8'b1111111;
DRAM[24491] = 8'b10000001;
DRAM[24492] = 8'b10000111;
DRAM[24493] = 8'b10001111;
DRAM[24494] = 8'b10011101;
DRAM[24495] = 8'b10101011;
DRAM[24496] = 8'b10111110;
DRAM[24497] = 8'b11010010;
DRAM[24498] = 8'b11011101;
DRAM[24499] = 8'b11100001;
DRAM[24500] = 8'b11101000;
DRAM[24501] = 8'b11100111;
DRAM[24502] = 8'b11100010;
DRAM[24503] = 8'b11100101;
DRAM[24504] = 8'b11110000;
DRAM[24505] = 8'b11100101;
DRAM[24506] = 8'b11011101;
DRAM[24507] = 8'b11010010;
DRAM[24508] = 8'b11000100;
DRAM[24509] = 8'b11000111;
DRAM[24510] = 8'b11001010;
DRAM[24511] = 8'b11000010;
DRAM[24512] = 8'b10011010;
DRAM[24513] = 8'b10010010;
DRAM[24514] = 8'b1101111;
DRAM[24515] = 8'b1010000;
DRAM[24516] = 8'b1001011;
DRAM[24517] = 8'b10001011;
DRAM[24518] = 8'b10010010;
DRAM[24519] = 8'b10010111;
DRAM[24520] = 8'b10100000;
DRAM[24521] = 8'b10101010;
DRAM[24522] = 8'b10111101;
DRAM[24523] = 8'b11101001;
DRAM[24524] = 8'b11110011;
DRAM[24525] = 8'b11110011;
DRAM[24526] = 8'b11111111;
DRAM[24527] = 8'b11100010;
DRAM[24528] = 8'b11010111;
DRAM[24529] = 8'b11101110;
DRAM[24530] = 8'b11100001;
DRAM[24531] = 8'b11011100;
DRAM[24532] = 8'b10101101;
DRAM[24533] = 8'b11001011;
DRAM[24534] = 8'b11000001;
DRAM[24535] = 8'b10111101;
DRAM[24536] = 8'b10100000;
DRAM[24537] = 8'b10111100;
DRAM[24538] = 8'b10110110;
DRAM[24539] = 8'b10011000;
DRAM[24540] = 8'b10111101;
DRAM[24541] = 8'b10100111;
DRAM[24542] = 8'b10011111;
DRAM[24543] = 8'b10111001;
DRAM[24544] = 8'b10110010;
DRAM[24545] = 8'b10001011;
DRAM[24546] = 8'b10111010;
DRAM[24547] = 8'b10010110;
DRAM[24548] = 8'b10011100;
DRAM[24549] = 8'b11001101;
DRAM[24550] = 8'b11011000;
DRAM[24551] = 8'b11001100;
DRAM[24552] = 8'b11101010;
DRAM[24553] = 8'b11100100;
DRAM[24554] = 8'b11000000;
DRAM[24555] = 8'b10011010;
DRAM[24556] = 8'b10001010;
DRAM[24557] = 8'b1110111;
DRAM[24558] = 8'b1101001;
DRAM[24559] = 8'b1110101;
DRAM[24560] = 8'b1101100;
DRAM[24561] = 8'b1101100;
DRAM[24562] = 8'b1101100;
DRAM[24563] = 8'b1101011;
DRAM[24564] = 8'b1101011;
DRAM[24565] = 8'b1101010;
DRAM[24566] = 8'b1101010;
DRAM[24567] = 8'b1101010;
DRAM[24568] = 8'b1101011;
DRAM[24569] = 8'b1101011;
DRAM[24570] = 8'b1101010;
DRAM[24571] = 8'b1101010;
DRAM[24572] = 8'b1101001;
DRAM[24573] = 8'b1101000;
DRAM[24574] = 8'b1100111;
DRAM[24575] = 8'b1100111;
DRAM[24576] = 8'b1111100;
DRAM[24577] = 8'b1111100;
DRAM[24578] = 8'b1111100;
DRAM[24579] = 8'b1111101;
DRAM[24580] = 8'b1111101;
DRAM[24581] = 8'b1111101;
DRAM[24582] = 8'b1111110;
DRAM[24583] = 8'b1111110;
DRAM[24584] = 8'b10000001;
DRAM[24585] = 8'b10000001;
DRAM[24586] = 8'b10000001;
DRAM[24587] = 8'b10000001;
DRAM[24588] = 8'b10000001;
DRAM[24589] = 8'b10000001;
DRAM[24590] = 8'b10000001;
DRAM[24591] = 8'b10000001;
DRAM[24592] = 8'b10000001;
DRAM[24593] = 8'b10000010;
DRAM[24594] = 8'b10000011;
DRAM[24595] = 8'b10000100;
DRAM[24596] = 8'b10000101;
DRAM[24597] = 8'b10000101;
DRAM[24598] = 8'b10000101;
DRAM[24599] = 8'b10000101;
DRAM[24600] = 8'b10001111;
DRAM[24601] = 8'b10010000;
DRAM[24602] = 8'b10010110;
DRAM[24603] = 8'b10111101;
DRAM[24604] = 8'b11001101;
DRAM[24605] = 8'b11110000;
DRAM[24606] = 8'b11100110;
DRAM[24607] = 8'b11010110;
DRAM[24608] = 8'b11011010;
DRAM[24609] = 8'b11010100;
DRAM[24610] = 8'b10100100;
DRAM[24611] = 8'b10101111;
DRAM[24612] = 8'b11010000;
DRAM[24613] = 8'b11000101;
DRAM[24614] = 8'b10111111;
DRAM[24615] = 8'b10111101;
DRAM[24616] = 8'b10100100;
DRAM[24617] = 8'b11000100;
DRAM[24618] = 8'b10111100;
DRAM[24619] = 8'b11000010;
DRAM[24620] = 8'b11011101;
DRAM[24621] = 8'b10101000;
DRAM[24622] = 8'b10111010;
DRAM[24623] = 8'b11100110;
DRAM[24624] = 8'b10110010;
DRAM[24625] = 8'b10110011;
DRAM[24626] = 8'b11011111;
DRAM[24627] = 8'b11001111;
DRAM[24628] = 8'b11000111;
DRAM[24629] = 8'b10111010;
DRAM[24630] = 8'b10111001;
DRAM[24631] = 8'b11000110;
DRAM[24632] = 8'b11010111;
DRAM[24633] = 8'b11000101;
DRAM[24634] = 8'b11011011;
DRAM[24635] = 8'b11100001;
DRAM[24636] = 8'b11000011;
DRAM[24637] = 8'b11001011;
DRAM[24638] = 8'b11101101;
DRAM[24639] = 8'b11101100;
DRAM[24640] = 8'b11101000;
DRAM[24641] = 8'b11010111;
DRAM[24642] = 8'b11011001;
DRAM[24643] = 8'b11100101;
DRAM[24644] = 8'b11010010;
DRAM[24645] = 8'b11100101;
DRAM[24646] = 8'b11001010;
DRAM[24647] = 8'b10111011;
DRAM[24648] = 8'b11000111;
DRAM[24649] = 8'b10011100;
DRAM[24650] = 8'b10110010;
DRAM[24651] = 8'b1110000;
DRAM[24652] = 8'b1010111;
DRAM[24653] = 8'b1101011;
DRAM[24654] = 8'b1110001;
DRAM[24655] = 8'b10000111;
DRAM[24656] = 8'b10001000;
DRAM[24657] = 8'b10001001;
DRAM[24658] = 8'b10010100;
DRAM[24659] = 8'b10100101;
DRAM[24660] = 8'b10101101;
DRAM[24661] = 8'b10101110;
DRAM[24662] = 8'b10110111;
DRAM[24663] = 8'b11000011;
DRAM[24664] = 8'b11000001;
DRAM[24665] = 8'b11001010;
DRAM[24666] = 8'b11001100;
DRAM[24667] = 8'b11000110;
DRAM[24668] = 8'b11000101;
DRAM[24669] = 8'b11001001;
DRAM[24670] = 8'b11000111;
DRAM[24671] = 8'b10111111;
DRAM[24672] = 8'b11000111;
DRAM[24673] = 8'b11000110;
DRAM[24674] = 8'b11001010;
DRAM[24675] = 8'b11001111;
DRAM[24676] = 8'b11001101;
DRAM[24677] = 8'b11000101;
DRAM[24678] = 8'b11000011;
DRAM[24679] = 8'b11000110;
DRAM[24680] = 8'b11001111;
DRAM[24681] = 8'b11001101;
DRAM[24682] = 8'b11000011;
DRAM[24683] = 8'b10111111;
DRAM[24684] = 8'b11000010;
DRAM[24685] = 8'b10111010;
DRAM[24686] = 8'b10110100;
DRAM[24687] = 8'b10111010;
DRAM[24688] = 8'b10110001;
DRAM[24689] = 8'b10011010;
DRAM[24690] = 8'b10101001;
DRAM[24691] = 8'b10010100;
DRAM[24692] = 8'b10011111;
DRAM[24693] = 8'b10001101;
DRAM[24694] = 8'b10110110;
DRAM[24695] = 8'b11000000;
DRAM[24696] = 8'b10110100;
DRAM[24697] = 8'b11000001;
DRAM[24698] = 8'b10111001;
DRAM[24699] = 8'b10010110;
DRAM[24700] = 8'b10100110;
DRAM[24701] = 8'b10110110;
DRAM[24702] = 8'b10011010;
DRAM[24703] = 8'b10100100;
DRAM[24704] = 8'b10010010;
DRAM[24705] = 8'b10011101;
DRAM[24706] = 8'b10100000;
DRAM[24707] = 8'b10011001;
DRAM[24708] = 8'b10011101;
DRAM[24709] = 8'b10101000;
DRAM[24710] = 8'b10100101;
DRAM[24711] = 8'b10011000;
DRAM[24712] = 8'b10101100;
DRAM[24713] = 8'b10100011;
DRAM[24714] = 8'b10101000;
DRAM[24715] = 8'b10011011;
DRAM[24716] = 8'b10101110;
DRAM[24717] = 8'b10100110;
DRAM[24718] = 8'b10101110;
DRAM[24719] = 8'b10100100;
DRAM[24720] = 8'b10100100;
DRAM[24721] = 8'b10101111;
DRAM[24722] = 8'b10011000;
DRAM[24723] = 8'b10011111;
DRAM[24724] = 8'b10101001;
DRAM[24725] = 8'b10011111;
DRAM[24726] = 8'b10100011;
DRAM[24727] = 8'b10010111;
DRAM[24728] = 8'b10011011;
DRAM[24729] = 8'b10011110;
DRAM[24730] = 8'b10011101;
DRAM[24731] = 8'b10010111;
DRAM[24732] = 8'b10010000;
DRAM[24733] = 8'b10001000;
DRAM[24734] = 8'b1111100;
DRAM[24735] = 8'b1110000;
DRAM[24736] = 8'b1101001;
DRAM[24737] = 8'b1110010;
DRAM[24738] = 8'b1101110;
DRAM[24739] = 8'b10000011;
DRAM[24740] = 8'b10000001;
DRAM[24741] = 8'b10010110;
DRAM[24742] = 8'b10001100;
DRAM[24743] = 8'b10001101;
DRAM[24744] = 8'b1110001;
DRAM[24745] = 8'b1110100;
DRAM[24746] = 8'b1110111;
DRAM[24747] = 8'b10000100;
DRAM[24748] = 8'b10010011;
DRAM[24749] = 8'b10011000;
DRAM[24750] = 8'b10100011;
DRAM[24751] = 8'b10111010;
DRAM[24752] = 8'b10101100;
DRAM[24753] = 8'b10110000;
DRAM[24754] = 8'b11000011;
DRAM[24755] = 8'b11100000;
DRAM[24756] = 8'b11110001;
DRAM[24757] = 8'b11101111;
DRAM[24758] = 8'b11101000;
DRAM[24759] = 8'b11100110;
DRAM[24760] = 8'b11100100;
DRAM[24761] = 8'b11110001;
DRAM[24762] = 8'b11101101;
DRAM[24763] = 8'b11011100;
DRAM[24764] = 8'b11001010;
DRAM[24765] = 8'b10110010;
DRAM[24766] = 8'b10011101;
DRAM[24767] = 8'b10011000;
DRAM[24768] = 8'b10010000;
DRAM[24769] = 8'b1110110;
DRAM[24770] = 8'b1110001;
DRAM[24771] = 8'b1100010;
DRAM[24772] = 8'b1010001;
DRAM[24773] = 8'b1101100;
DRAM[24774] = 8'b10010011;
DRAM[24775] = 8'b10101011;
DRAM[24776] = 8'b10111001;
DRAM[24777] = 8'b10011100;
DRAM[24778] = 8'b10111010;
DRAM[24779] = 8'b11011010;
DRAM[24780] = 8'b11101111;
DRAM[24781] = 8'b11111001;
DRAM[24782] = 8'b11101100;
DRAM[24783] = 8'b11110101;
DRAM[24784] = 8'b11010101;
DRAM[24785] = 8'b11100111;
DRAM[24786] = 8'b11011000;
DRAM[24787] = 8'b11100000;
DRAM[24788] = 8'b10110111;
DRAM[24789] = 8'b10111001;
DRAM[24790] = 8'b11001101;
DRAM[24791] = 8'b10111111;
DRAM[24792] = 8'b10100011;
DRAM[24793] = 8'b10100110;
DRAM[24794] = 8'b11000010;
DRAM[24795] = 8'b10110000;
DRAM[24796] = 8'b10100011;
DRAM[24797] = 8'b10110101;
DRAM[24798] = 8'b10101001;
DRAM[24799] = 8'b10100101;
DRAM[24800] = 8'b10110101;
DRAM[24801] = 8'b10011101;
DRAM[24802] = 8'b10100100;
DRAM[24803] = 8'b10100000;
DRAM[24804] = 8'b10100110;
DRAM[24805] = 8'b10111001;
DRAM[24806] = 8'b11000010;
DRAM[24807] = 8'b11100100;
DRAM[24808] = 8'b11100010;
DRAM[24809] = 8'b11100000;
DRAM[24810] = 8'b10110001;
DRAM[24811] = 8'b10011010;
DRAM[24812] = 8'b10001011;
DRAM[24813] = 8'b1110101;
DRAM[24814] = 8'b1110110;
DRAM[24815] = 8'b1101011;
DRAM[24816] = 8'b1101101;
DRAM[24817] = 8'b1101101;
DRAM[24818] = 8'b1101100;
DRAM[24819] = 8'b1101100;
DRAM[24820] = 8'b1101100;
DRAM[24821] = 8'b1101011;
DRAM[24822] = 8'b1101011;
DRAM[24823] = 8'b1101011;
DRAM[24824] = 8'b1101010;
DRAM[24825] = 8'b1101010;
DRAM[24826] = 8'b1101001;
DRAM[24827] = 8'b1101001;
DRAM[24828] = 8'b1101001;
DRAM[24829] = 8'b1101000;
DRAM[24830] = 8'b1101000;
DRAM[24831] = 8'b1101000;
DRAM[24832] = 8'b1111100;
DRAM[24833] = 8'b1111100;
DRAM[24834] = 8'b1111101;
DRAM[24835] = 8'b1111101;
DRAM[24836] = 8'b1111101;
DRAM[24837] = 8'b1111110;
DRAM[24838] = 8'b1111110;
DRAM[24839] = 8'b1111110;
DRAM[24840] = 8'b10000001;
DRAM[24841] = 8'b10000001;
DRAM[24842] = 8'b10000001;
DRAM[24843] = 8'b10000001;
DRAM[24844] = 8'b10000001;
DRAM[24845] = 8'b10000010;
DRAM[24846] = 8'b10000010;
DRAM[24847] = 8'b10000010;
DRAM[24848] = 8'b10000010;
DRAM[24849] = 8'b10000011;
DRAM[24850] = 8'b10000100;
DRAM[24851] = 8'b10000101;
DRAM[24852] = 8'b10000110;
DRAM[24853] = 8'b10000110;
DRAM[24854] = 8'b10000110;
DRAM[24855] = 8'b10000110;
DRAM[24856] = 8'b10000110;
DRAM[24857] = 8'b10010010;
DRAM[24858] = 8'b10110000;
DRAM[24859] = 8'b10011011;
DRAM[24860] = 8'b11000001;
DRAM[24861] = 8'b11010101;
DRAM[24862] = 8'b11110101;
DRAM[24863] = 8'b11011100;
DRAM[24864] = 8'b11011001;
DRAM[24865] = 8'b11000000;
DRAM[24866] = 8'b10111001;
DRAM[24867] = 8'b11001111;
DRAM[24868] = 8'b10111110;
DRAM[24869] = 8'b10101111;
DRAM[24870] = 8'b11000010;
DRAM[24871] = 8'b10110011;
DRAM[24872] = 8'b10100011;
DRAM[24873] = 8'b11001001;
DRAM[24874] = 8'b11000100;
DRAM[24875] = 8'b10110111;
DRAM[24876] = 8'b10110100;
DRAM[24877] = 8'b10111111;
DRAM[24878] = 8'b11000110;
DRAM[24879] = 8'b11000001;
DRAM[24880] = 8'b10110001;
DRAM[24881] = 8'b11000000;
DRAM[24882] = 8'b11010011;
DRAM[24883] = 8'b10110111;
DRAM[24884] = 8'b11000111;
DRAM[24885] = 8'b10111110;
DRAM[24886] = 8'b10110011;
DRAM[24887] = 8'b11000110;
DRAM[24888] = 8'b11010100;
DRAM[24889] = 8'b11001011;
DRAM[24890] = 8'b11011111;
DRAM[24891] = 8'b11011100;
DRAM[24892] = 8'b11001110;
DRAM[24893] = 8'b11010010;
DRAM[24894] = 8'b11101110;
DRAM[24895] = 8'b11101011;
DRAM[24896] = 8'b11100100;
DRAM[24897] = 8'b11011010;
DRAM[24898] = 8'b11011010;
DRAM[24899] = 8'b11100010;
DRAM[24900] = 8'b11010111;
DRAM[24901] = 8'b11100101;
DRAM[24902] = 8'b11000101;
DRAM[24903] = 8'b10111000;
DRAM[24904] = 8'b11010110;
DRAM[24905] = 8'b10101010;
DRAM[24906] = 8'b10110010;
DRAM[24907] = 8'b1101000;
DRAM[24908] = 8'b1010000;
DRAM[24909] = 8'b1101000;
DRAM[24910] = 8'b1101110;
DRAM[24911] = 8'b1111111;
DRAM[24912] = 8'b10000100;
DRAM[24913] = 8'b10001010;
DRAM[24914] = 8'b10010111;
DRAM[24915] = 8'b10100101;
DRAM[24916] = 8'b10101110;
DRAM[24917] = 8'b10110100;
DRAM[24918] = 8'b10111110;
DRAM[24919] = 8'b11000111;
DRAM[24920] = 8'b10111010;
DRAM[24921] = 8'b10111101;
DRAM[24922] = 8'b10111111;
DRAM[24923] = 8'b10111111;
DRAM[24924] = 8'b11000000;
DRAM[24925] = 8'b11000001;
DRAM[24926] = 8'b10111110;
DRAM[24927] = 8'b10111000;
DRAM[24928] = 8'b10110011;
DRAM[24929] = 8'b10111001;
DRAM[24930] = 8'b11000111;
DRAM[24931] = 8'b11010111;
DRAM[24932] = 8'b11011101;
DRAM[24933] = 8'b11010111;
DRAM[24934] = 8'b11010000;
DRAM[24935] = 8'b11001110;
DRAM[24936] = 8'b11001010;
DRAM[24937] = 8'b11001010;
DRAM[24938] = 8'b11000010;
DRAM[24939] = 8'b11000000;
DRAM[24940] = 8'b11000100;
DRAM[24941] = 8'b10111100;
DRAM[24942] = 8'b10110101;
DRAM[24943] = 8'b10111011;
DRAM[24944] = 8'b11000001;
DRAM[24945] = 8'b10011001;
DRAM[24946] = 8'b10101111;
DRAM[24947] = 8'b10110011;
DRAM[24948] = 8'b10010111;
DRAM[24949] = 8'b10010100;
DRAM[24950] = 8'b10110101;
DRAM[24951] = 8'b10100001;
DRAM[24952] = 8'b10101101;
DRAM[24953] = 8'b10110011;
DRAM[24954] = 8'b10110110;
DRAM[24955] = 8'b10100001;
DRAM[24956] = 8'b10100101;
DRAM[24957] = 8'b10101000;
DRAM[24958] = 8'b10010101;
DRAM[24959] = 8'b10100011;
DRAM[24960] = 8'b10010011;
DRAM[24961] = 8'b10010110;
DRAM[24962] = 8'b10011000;
DRAM[24963] = 8'b10011001;
DRAM[24964] = 8'b10011010;
DRAM[24965] = 8'b10011110;
DRAM[24966] = 8'b10100010;
DRAM[24967] = 8'b10100011;
DRAM[24968] = 8'b10101010;
DRAM[24969] = 8'b10100101;
DRAM[24970] = 8'b10101101;
DRAM[24971] = 8'b10100010;
DRAM[24972] = 8'b10101111;
DRAM[24973] = 8'b10100110;
DRAM[24974] = 8'b10101100;
DRAM[24975] = 8'b10100101;
DRAM[24976] = 8'b10011000;
DRAM[24977] = 8'b10100100;
DRAM[24978] = 8'b10011000;
DRAM[24979] = 8'b10100001;
DRAM[24980] = 8'b10011111;
DRAM[24981] = 8'b10001011;
DRAM[24982] = 8'b10011001;
DRAM[24983] = 8'b10100101;
DRAM[24984] = 8'b10010111;
DRAM[24985] = 8'b10011101;
DRAM[24986] = 8'b10010111;
DRAM[24987] = 8'b10001001;
DRAM[24988] = 8'b10000110;
DRAM[24989] = 8'b10001010;
DRAM[24990] = 8'b1111100;
DRAM[24991] = 8'b1100101;
DRAM[24992] = 8'b1110000;
DRAM[24993] = 8'b1100110;
DRAM[24994] = 8'b1011000;
DRAM[24995] = 8'b1110010;
DRAM[24996] = 8'b1111011;
DRAM[24997] = 8'b10001000;
DRAM[24998] = 8'b1101111;
DRAM[24999] = 8'b1100010;
DRAM[25000] = 8'b1000111;
DRAM[25001] = 8'b1101010;
DRAM[25002] = 8'b1111111;
DRAM[25003] = 8'b10000010;
DRAM[25004] = 8'b10001100;
DRAM[25005] = 8'b10011000;
DRAM[25006] = 8'b10100000;
DRAM[25007] = 8'b10100111;
DRAM[25008] = 8'b10111100;
DRAM[25009] = 8'b11000101;
DRAM[25010] = 8'b11001010;
DRAM[25011] = 8'b11000110;
DRAM[25012] = 8'b11000101;
DRAM[25013] = 8'b11010010;
DRAM[25014] = 8'b11101001;
DRAM[25015] = 8'b11111010;
DRAM[25016] = 8'b11100000;
DRAM[25017] = 8'b11101011;
DRAM[25018] = 8'b11100111;
DRAM[25019] = 8'b11011100;
DRAM[25020] = 8'b11010101;
DRAM[25021] = 8'b11001001;
DRAM[25022] = 8'b10111101;
DRAM[25023] = 8'b10111101;
DRAM[25024] = 8'b10100111;
DRAM[25025] = 8'b10001100;
DRAM[25026] = 8'b1111100;
DRAM[25027] = 8'b1100001;
DRAM[25028] = 8'b1001010;
DRAM[25029] = 8'b1011111;
DRAM[25030] = 8'b10000101;
DRAM[25031] = 8'b10010101;
DRAM[25032] = 8'b10110011;
DRAM[25033] = 8'b10011110;
DRAM[25034] = 8'b10111011;
DRAM[25035] = 8'b11011011;
DRAM[25036] = 8'b11101111;
DRAM[25037] = 8'b11110111;
DRAM[25038] = 8'b11101001;
DRAM[25039] = 8'b11110010;
DRAM[25040] = 8'b11011111;
DRAM[25041] = 8'b11011100;
DRAM[25042] = 8'b11100001;
DRAM[25043] = 8'b11010111;
DRAM[25044] = 8'b11001000;
DRAM[25045] = 8'b10110000;
DRAM[25046] = 8'b11000010;
DRAM[25047] = 8'b10111101;
DRAM[25048] = 8'b10100100;
DRAM[25049] = 8'b10101001;
DRAM[25050] = 8'b10111001;
DRAM[25051] = 8'b10101111;
DRAM[25052] = 8'b10100110;
DRAM[25053] = 8'b10101110;
DRAM[25054] = 8'b10101101;
DRAM[25055] = 8'b10101010;
DRAM[25056] = 8'b10101000;
DRAM[25057] = 8'b10010110;
DRAM[25058] = 8'b10011111;
DRAM[25059] = 8'b10011110;
DRAM[25060] = 8'b10100111;
DRAM[25061] = 8'b10111010;
DRAM[25062] = 8'b11000100;
DRAM[25063] = 8'b11100011;
DRAM[25064] = 8'b11010110;
DRAM[25065] = 8'b11100000;
DRAM[25066] = 8'b10111001;
DRAM[25067] = 8'b10010111;
DRAM[25068] = 8'b10000000;
DRAM[25069] = 8'b1110001;
DRAM[25070] = 8'b1110101;
DRAM[25071] = 8'b1101000;
DRAM[25072] = 8'b1101101;
DRAM[25073] = 8'b1101101;
DRAM[25074] = 8'b1101101;
DRAM[25075] = 8'b1101100;
DRAM[25076] = 8'b1101100;
DRAM[25077] = 8'b1101100;
DRAM[25078] = 8'b1101011;
DRAM[25079] = 8'b1101011;
DRAM[25080] = 8'b1101010;
DRAM[25081] = 8'b1101010;
DRAM[25082] = 8'b1101010;
DRAM[25083] = 8'b1101001;
DRAM[25084] = 8'b1101001;
DRAM[25085] = 8'b1101001;
DRAM[25086] = 8'b1101000;
DRAM[25087] = 8'b1101000;
DRAM[25088] = 8'b1111101;
DRAM[25089] = 8'b1111101;
DRAM[25090] = 8'b1111101;
DRAM[25091] = 8'b1111110;
DRAM[25092] = 8'b1111110;
DRAM[25093] = 8'b1111110;
DRAM[25094] = 8'b1111111;
DRAM[25095] = 8'b1111111;
DRAM[25096] = 8'b10000000;
DRAM[25097] = 8'b10000001;
DRAM[25098] = 8'b10000001;
DRAM[25099] = 8'b10000010;
DRAM[25100] = 8'b10000010;
DRAM[25101] = 8'b10000011;
DRAM[25102] = 8'b10000011;
DRAM[25103] = 8'b10000011;
DRAM[25104] = 8'b10000100;
DRAM[25105] = 8'b10000100;
DRAM[25106] = 8'b10000101;
DRAM[25107] = 8'b10000110;
DRAM[25108] = 8'b10000110;
DRAM[25109] = 8'b10000111;
DRAM[25110] = 8'b10001000;
DRAM[25111] = 8'b10001000;
DRAM[25112] = 8'b10001100;
DRAM[25113] = 8'b10011000;
DRAM[25114] = 8'b10010110;
DRAM[25115] = 8'b10011100;
DRAM[25116] = 8'b10110101;
DRAM[25117] = 8'b11100011;
DRAM[25118] = 8'b11101011;
DRAM[25119] = 8'b11011100;
DRAM[25120] = 8'b11010001;
DRAM[25121] = 8'b11000001;
DRAM[25122] = 8'b10111001;
DRAM[25123] = 8'b10111110;
DRAM[25124] = 8'b10110010;
DRAM[25125] = 8'b10110111;
DRAM[25126] = 8'b11000000;
DRAM[25127] = 8'b10011100;
DRAM[25128] = 8'b11000100;
DRAM[25129] = 8'b10111111;
DRAM[25130] = 8'b10111010;
DRAM[25131] = 8'b10110110;
DRAM[25132] = 8'b10011101;
DRAM[25133] = 8'b11000111;
DRAM[25134] = 8'b11001000;
DRAM[25135] = 8'b11000100;
DRAM[25136] = 8'b10101100;
DRAM[25137] = 8'b11000001;
DRAM[25138] = 8'b10111111;
DRAM[25139] = 8'b10011110;
DRAM[25140] = 8'b11000001;
DRAM[25141] = 8'b10111100;
DRAM[25142] = 8'b10110001;
DRAM[25143] = 8'b11000111;
DRAM[25144] = 8'b11000100;
DRAM[25145] = 8'b11001001;
DRAM[25146] = 8'b11011010;
DRAM[25147] = 8'b11001100;
DRAM[25148] = 8'b11011000;
DRAM[25149] = 8'b11010111;
DRAM[25150] = 8'b11101011;
DRAM[25151] = 8'b11100111;
DRAM[25152] = 8'b11100001;
DRAM[25153] = 8'b11011111;
DRAM[25154] = 8'b11011100;
DRAM[25155] = 8'b11011100;
DRAM[25156] = 8'b11011111;
DRAM[25157] = 8'b11100111;
DRAM[25158] = 8'b11000010;
DRAM[25159] = 8'b10111010;
DRAM[25160] = 8'b10111110;
DRAM[25161] = 8'b10011111;
DRAM[25162] = 8'b10100110;
DRAM[25163] = 8'b1100000;
DRAM[25164] = 8'b1010011;
DRAM[25165] = 8'b1110001;
DRAM[25166] = 8'b1111001;
DRAM[25167] = 8'b10000011;
DRAM[25168] = 8'b10010000;
DRAM[25169] = 8'b10011011;
DRAM[25170] = 8'b10100110;
DRAM[25171] = 8'b10101100;
DRAM[25172] = 8'b10110010;
DRAM[25173] = 8'b10111010;
DRAM[25174] = 8'b11000001;
DRAM[25175] = 8'b11000011;
DRAM[25176] = 8'b11010100;
DRAM[25177] = 8'b11001110;
DRAM[25178] = 8'b11001011;
DRAM[25179] = 8'b11001101;
DRAM[25180] = 8'b11001100;
DRAM[25181] = 8'b11000110;
DRAM[25182] = 8'b11000000;
DRAM[25183] = 8'b10111110;
DRAM[25184] = 8'b11010011;
DRAM[25185] = 8'b11010000;
DRAM[25186] = 8'b11010001;
DRAM[25187] = 8'b11011000;
DRAM[25188] = 8'b11011100;
DRAM[25189] = 8'b11011010;
DRAM[25190] = 8'b11010110;
DRAM[25191] = 8'b11010101;
DRAM[25192] = 8'b11000110;
DRAM[25193] = 8'b11000101;
DRAM[25194] = 8'b10111100;
DRAM[25195] = 8'b10111000;
DRAM[25196] = 8'b10111001;
DRAM[25197] = 8'b10101101;
DRAM[25198] = 8'b10100011;
DRAM[25199] = 8'b10100111;
DRAM[25200] = 8'b10110111;
DRAM[25201] = 8'b10011111;
DRAM[25202] = 8'b10100101;
DRAM[25203] = 8'b10110010;
DRAM[25204] = 8'b10011001;
DRAM[25205] = 8'b10011101;
DRAM[25206] = 8'b10100101;
DRAM[25207] = 8'b10011010;
DRAM[25208] = 8'b10110001;
DRAM[25209] = 8'b10110001;
DRAM[25210] = 8'b10111101;
DRAM[25211] = 8'b10110101;
DRAM[25212] = 8'b10101010;
DRAM[25213] = 8'b10100101;
DRAM[25214] = 8'b10011111;
DRAM[25215] = 8'b10101110;
DRAM[25216] = 8'b10010001;
DRAM[25217] = 8'b10001111;
DRAM[25218] = 8'b10010011;
DRAM[25219] = 8'b10011000;
DRAM[25220] = 8'b10010110;
DRAM[25221] = 8'b10010100;
DRAM[25222] = 8'b10011110;
DRAM[25223] = 8'b10101101;
DRAM[25224] = 8'b10100010;
DRAM[25225] = 8'b10100011;
DRAM[25226] = 8'b10101100;
DRAM[25227] = 8'b10100110;
DRAM[25228] = 8'b10101011;
DRAM[25229] = 8'b10011111;
DRAM[25230] = 8'b10100011;
DRAM[25231] = 8'b10100000;
DRAM[25232] = 8'b10011101;
DRAM[25233] = 8'b10011110;
DRAM[25234] = 8'b10010110;
DRAM[25235] = 8'b10100011;
DRAM[25236] = 8'b10100000;
DRAM[25237] = 8'b10000111;
DRAM[25238] = 8'b10010010;
DRAM[25239] = 8'b10101010;
DRAM[25240] = 8'b10011100;
DRAM[25241] = 8'b10100100;
DRAM[25242] = 8'b10011011;
DRAM[25243] = 8'b10001000;
DRAM[25244] = 8'b10001010;
DRAM[25245] = 8'b10011000;
DRAM[25246] = 8'b10001100;
DRAM[25247] = 8'b1101110;
DRAM[25248] = 8'b1111000;
DRAM[25249] = 8'b1100100;
DRAM[25250] = 8'b1010111;
DRAM[25251] = 8'b1110000;
DRAM[25252] = 8'b1111000;
DRAM[25253] = 8'b1110100;
DRAM[25254] = 8'b1010110;
DRAM[25255] = 8'b1001001;
DRAM[25256] = 8'b1110011;
DRAM[25257] = 8'b10000001;
DRAM[25258] = 8'b10000010;
DRAM[25259] = 8'b10000100;
DRAM[25260] = 8'b10011010;
DRAM[25261] = 8'b10101010;
DRAM[25262] = 8'b10100111;
DRAM[25263] = 8'b10100010;
DRAM[25264] = 8'b10101010;
DRAM[25265] = 8'b10110111;
DRAM[25266] = 8'b10111110;
DRAM[25267] = 8'b10111111;
DRAM[25268] = 8'b11001010;
DRAM[25269] = 8'b11011110;
DRAM[25270] = 8'b11101000;
DRAM[25271] = 8'b11100110;
DRAM[25272] = 8'b11110001;
DRAM[25273] = 8'b11111001;
DRAM[25274] = 8'b11110010;
DRAM[25275] = 8'b11100101;
DRAM[25276] = 8'b11100000;
DRAM[25277] = 8'b11010011;
DRAM[25278] = 8'b11000011;
DRAM[25279] = 8'b10111110;
DRAM[25280] = 8'b10110010;
DRAM[25281] = 8'b10011110;
DRAM[25282] = 8'b10001011;
DRAM[25283] = 8'b1110000;
DRAM[25284] = 8'b1010111;
DRAM[25285] = 8'b1101011;
DRAM[25286] = 8'b10001111;
DRAM[25287] = 8'b10010101;
DRAM[25288] = 8'b10101011;
DRAM[25289] = 8'b10100010;
DRAM[25290] = 8'b10111100;
DRAM[25291] = 8'b11011011;
DRAM[25292] = 8'b11110000;
DRAM[25293] = 8'b11110010;
DRAM[25294] = 8'b11100101;
DRAM[25295] = 8'b11101100;
DRAM[25296] = 8'b11101011;
DRAM[25297] = 8'b11010100;
DRAM[25298] = 8'b11101100;
DRAM[25299] = 8'b11001101;
DRAM[25300] = 8'b11011011;
DRAM[25301] = 8'b10110001;
DRAM[25302] = 8'b10111000;
DRAM[25303] = 8'b10110111;
DRAM[25304] = 8'b10100110;
DRAM[25305] = 8'b10101101;
DRAM[25306] = 8'b10101001;
DRAM[25307] = 8'b10101100;
DRAM[25308] = 8'b10100110;
DRAM[25309] = 8'b10100001;
DRAM[25310] = 8'b10101100;
DRAM[25311] = 8'b10101101;
DRAM[25312] = 8'b10011100;
DRAM[25313] = 8'b10010010;
DRAM[25314] = 8'b10011010;
DRAM[25315] = 8'b10011101;
DRAM[25316] = 8'b10100110;
DRAM[25317] = 8'b10111000;
DRAM[25318] = 8'b11000100;
DRAM[25319] = 8'b11011101;
DRAM[25320] = 8'b11000010;
DRAM[25321] = 8'b11010001;
DRAM[25322] = 8'b10111010;
DRAM[25323] = 8'b10010101;
DRAM[25324] = 8'b1111000;
DRAM[25325] = 8'b1101111;
DRAM[25326] = 8'b1110111;
DRAM[25327] = 8'b1101011;
DRAM[25328] = 8'b1101110;
DRAM[25329] = 8'b1101110;
DRAM[25330] = 8'b1101101;
DRAM[25331] = 8'b1101101;
DRAM[25332] = 8'b1101101;
DRAM[25333] = 8'b1101100;
DRAM[25334] = 8'b1101100;
DRAM[25335] = 8'b1101100;
DRAM[25336] = 8'b1101011;
DRAM[25337] = 8'b1101011;
DRAM[25338] = 8'b1101010;
DRAM[25339] = 8'b1101010;
DRAM[25340] = 8'b1101010;
DRAM[25341] = 8'b1101001;
DRAM[25342] = 8'b1101001;
DRAM[25343] = 8'b1101001;
DRAM[25344] = 8'b1111110;
DRAM[25345] = 8'b1111110;
DRAM[25346] = 8'b1111110;
DRAM[25347] = 8'b1111110;
DRAM[25348] = 8'b1111111;
DRAM[25349] = 8'b1111111;
DRAM[25350] = 8'b1111111;
DRAM[25351] = 8'b10000000;
DRAM[25352] = 8'b10000001;
DRAM[25353] = 8'b10000001;
DRAM[25354] = 8'b10000010;
DRAM[25355] = 8'b10000010;
DRAM[25356] = 8'b10000011;
DRAM[25357] = 8'b10000100;
DRAM[25358] = 8'b10000100;
DRAM[25359] = 8'b10000100;
DRAM[25360] = 8'b10000101;
DRAM[25361] = 8'b10000101;
DRAM[25362] = 8'b10000110;
DRAM[25363] = 8'b10000110;
DRAM[25364] = 8'b10000111;
DRAM[25365] = 8'b10001000;
DRAM[25366] = 8'b10001001;
DRAM[25367] = 8'b10001010;
DRAM[25368] = 8'b10010011;
DRAM[25369] = 8'b10010010;
DRAM[25370] = 8'b10000011;
DRAM[25371] = 8'b10101101;
DRAM[25372] = 8'b11000000;
DRAM[25373] = 8'b11100101;
DRAM[25374] = 8'b11011001;
DRAM[25375] = 8'b11100000;
DRAM[25376] = 8'b11010000;
DRAM[25377] = 8'b11001101;
DRAM[25378] = 8'b10101110;
DRAM[25379] = 8'b10101000;
DRAM[25380] = 8'b10111110;
DRAM[25381] = 8'b10110111;
DRAM[25382] = 8'b10101000;
DRAM[25383] = 8'b10101111;
DRAM[25384] = 8'b11000101;
DRAM[25385] = 8'b10110001;
DRAM[25386] = 8'b10111000;
DRAM[25387] = 8'b10110111;
DRAM[25388] = 8'b10101100;
DRAM[25389] = 8'b11001001;
DRAM[25390] = 8'b10111111;
DRAM[25391] = 8'b11000111;
DRAM[25392] = 8'b10101111;
DRAM[25393] = 8'b10110100;
DRAM[25394] = 8'b10110100;
DRAM[25395] = 8'b10100001;
DRAM[25396] = 8'b10111011;
DRAM[25397] = 8'b10110110;
DRAM[25398] = 8'b10111100;
DRAM[25399] = 8'b11001100;
DRAM[25400] = 8'b10110110;
DRAM[25401] = 8'b11000111;
DRAM[25402] = 8'b11010011;
DRAM[25403] = 8'b10111111;
DRAM[25404] = 8'b11011111;
DRAM[25405] = 8'b11011110;
DRAM[25406] = 8'b11101001;
DRAM[25407] = 8'b11100101;
DRAM[25408] = 8'b11100000;
DRAM[25409] = 8'b11100010;
DRAM[25410] = 8'b11011100;
DRAM[25411] = 8'b11010101;
DRAM[25412] = 8'b11100101;
DRAM[25413] = 8'b11101001;
DRAM[25414] = 8'b11000101;
DRAM[25415] = 8'b10111111;
DRAM[25416] = 8'b10111000;
DRAM[25417] = 8'b10101011;
DRAM[25418] = 8'b10110001;
DRAM[25419] = 8'b1101011;
DRAM[25420] = 8'b1011100;
DRAM[25421] = 8'b1101110;
DRAM[25422] = 8'b1101101;
DRAM[25423] = 8'b1101101;
DRAM[25424] = 8'b1111111;
DRAM[25425] = 8'b10010000;
DRAM[25426] = 8'b10100000;
DRAM[25427] = 8'b10101000;
DRAM[25428] = 8'b10110100;
DRAM[25429] = 8'b11000110;
DRAM[25430] = 8'b11010001;
DRAM[25431] = 8'b11010010;
DRAM[25432] = 8'b11011000;
DRAM[25433] = 8'b11001101;
DRAM[25434] = 8'b11001010;
DRAM[25435] = 8'b11010010;
DRAM[25436] = 8'b11010110;
DRAM[25437] = 8'b11010011;
DRAM[25438] = 8'b11010010;
DRAM[25439] = 8'b11010111;
DRAM[25440] = 8'b11110010;
DRAM[25441] = 8'b11101001;
DRAM[25442] = 8'b11011111;
DRAM[25443] = 8'b11011010;
DRAM[25444] = 8'b11011000;
DRAM[25445] = 8'b11010101;
DRAM[25446] = 8'b11001111;
DRAM[25447] = 8'b11001011;
DRAM[25448] = 8'b11001101;
DRAM[25449] = 8'b11001100;
DRAM[25450] = 8'b11000011;
DRAM[25451] = 8'b10111110;
DRAM[25452] = 8'b10111111;
DRAM[25453] = 8'b10110011;
DRAM[25454] = 8'b10101000;
DRAM[25455] = 8'b10101011;
DRAM[25456] = 8'b10110001;
DRAM[25457] = 8'b11000000;
DRAM[25458] = 8'b10101010;
DRAM[25459] = 8'b10011110;
DRAM[25460] = 8'b10110111;
DRAM[25461] = 8'b10101000;
DRAM[25462] = 8'b10011010;
DRAM[25463] = 8'b10110101;
DRAM[25464] = 8'b10100101;
DRAM[25465] = 8'b10100110;
DRAM[25466] = 8'b10110000;
DRAM[25467] = 8'b10101001;
DRAM[25468] = 8'b10011001;
DRAM[25469] = 8'b10011001;
DRAM[25470] = 8'b10100000;
DRAM[25471] = 8'b10100100;
DRAM[25472] = 8'b10001100;
DRAM[25473] = 8'b10010001;
DRAM[25474] = 8'b10010110;
DRAM[25475] = 8'b10010110;
DRAM[25476] = 8'b10010010;
DRAM[25477] = 8'b10010010;
DRAM[25478] = 8'b10011110;
DRAM[25479] = 8'b10101011;
DRAM[25480] = 8'b10011101;
DRAM[25481] = 8'b10100010;
DRAM[25482] = 8'b10101100;
DRAM[25483] = 8'b10101101;
DRAM[25484] = 8'b10101001;
DRAM[25485] = 8'b10011101;
DRAM[25486] = 8'b10011100;
DRAM[25487] = 8'b10011101;
DRAM[25488] = 8'b10101001;
DRAM[25489] = 8'b10011110;
DRAM[25490] = 8'b10010000;
DRAM[25491] = 8'b10011011;
DRAM[25492] = 8'b10100100;
DRAM[25493] = 8'b10010101;
DRAM[25494] = 8'b10001110;
DRAM[25495] = 8'b10010110;
DRAM[25496] = 8'b10010000;
DRAM[25497] = 8'b10010100;
DRAM[25498] = 8'b10001100;
DRAM[25499] = 8'b1111111;
DRAM[25500] = 8'b10000001;
DRAM[25501] = 8'b10001100;
DRAM[25502] = 8'b10000100;
DRAM[25503] = 8'b1110000;
DRAM[25504] = 8'b1110100;
DRAM[25505] = 8'b1100111;
DRAM[25506] = 8'b1100110;
DRAM[25507] = 8'b1111001;
DRAM[25508] = 8'b1110100;
DRAM[25509] = 8'b1011110;
DRAM[25510] = 8'b1001111;
DRAM[25511] = 8'b1010100;
DRAM[25512] = 8'b1111111;
DRAM[25513] = 8'b1110000;
DRAM[25514] = 8'b1100110;
DRAM[25515] = 8'b1111001;
DRAM[25516] = 8'b10010100;
DRAM[25517] = 8'b10011000;
DRAM[25518] = 8'b10010111;
DRAM[25519] = 8'b10100100;
DRAM[25520] = 8'b10100011;
DRAM[25521] = 8'b10101010;
DRAM[25522] = 8'b10110100;
DRAM[25523] = 8'b11000000;
DRAM[25524] = 8'b11001110;
DRAM[25525] = 8'b11010111;
DRAM[25526] = 8'b11010100;
DRAM[25527] = 8'b11001100;
DRAM[25528] = 8'b11100011;
DRAM[25529] = 8'b11101011;
DRAM[25530] = 8'b11100110;
DRAM[25531] = 8'b11011101;
DRAM[25532] = 8'b11010111;
DRAM[25533] = 8'b11000100;
DRAM[25534] = 8'b10101001;
DRAM[25535] = 8'b10011101;
DRAM[25536] = 8'b10011000;
DRAM[25537] = 8'b10001111;
DRAM[25538] = 8'b1111111;
DRAM[25539] = 8'b1101011;
DRAM[25540] = 8'b1010100;
DRAM[25541] = 8'b1100100;
DRAM[25542] = 8'b10001000;
DRAM[25543] = 8'b10000101;
DRAM[25544] = 8'b10100001;
DRAM[25545] = 8'b10100110;
DRAM[25546] = 8'b10111011;
DRAM[25547] = 8'b11011001;
DRAM[25548] = 8'b11110000;
DRAM[25549] = 8'b11101111;
DRAM[25550] = 8'b11100011;
DRAM[25551] = 8'b11101000;
DRAM[25552] = 8'b11110000;
DRAM[25553] = 8'b11010101;
DRAM[25554] = 8'b11101100;
DRAM[25555] = 8'b11001010;
DRAM[25556] = 8'b11011111;
DRAM[25557] = 8'b11000101;
DRAM[25558] = 8'b10110110;
DRAM[25559] = 8'b10101111;
DRAM[25560] = 8'b10101000;
DRAM[25561] = 8'b10110000;
DRAM[25562] = 8'b10011101;
DRAM[25563] = 8'b10100111;
DRAM[25564] = 8'b10100110;
DRAM[25565] = 8'b10010100;
DRAM[25566] = 8'b10100110;
DRAM[25567] = 8'b10101010;
DRAM[25568] = 8'b10011001;
DRAM[25569] = 8'b10010101;
DRAM[25570] = 8'b10011000;
DRAM[25571] = 8'b10011100;
DRAM[25572] = 8'b10100101;
DRAM[25573] = 8'b10110101;
DRAM[25574] = 8'b11000100;
DRAM[25575] = 8'b11010100;
DRAM[25576] = 8'b10101111;
DRAM[25577] = 8'b10110010;
DRAM[25578] = 8'b10101010;
DRAM[25579] = 8'b10010101;
DRAM[25580] = 8'b1111011;
DRAM[25581] = 8'b1110010;
DRAM[25582] = 8'b1110111;
DRAM[25583] = 8'b1110011;
DRAM[25584] = 8'b1101111;
DRAM[25585] = 8'b1101110;
DRAM[25586] = 8'b1101110;
DRAM[25587] = 8'b1101110;
DRAM[25588] = 8'b1101101;
DRAM[25589] = 8'b1101101;
DRAM[25590] = 8'b1101101;
DRAM[25591] = 8'b1101101;
DRAM[25592] = 8'b1101100;
DRAM[25593] = 8'b1101011;
DRAM[25594] = 8'b1101011;
DRAM[25595] = 8'b1101011;
DRAM[25596] = 8'b1101010;
DRAM[25597] = 8'b1101010;
DRAM[25598] = 8'b1101010;
DRAM[25599] = 8'b1101010;
DRAM[25600] = 8'b1111110;
DRAM[25601] = 8'b1111111;
DRAM[25602] = 8'b1111111;
DRAM[25603] = 8'b1111111;
DRAM[25604] = 8'b10000000;
DRAM[25605] = 8'b10000000;
DRAM[25606] = 8'b10000000;
DRAM[25607] = 8'b10000000;
DRAM[25608] = 8'b10000010;
DRAM[25609] = 8'b10000010;
DRAM[25610] = 8'b10000011;
DRAM[25611] = 8'b10000011;
DRAM[25612] = 8'b10000100;
DRAM[25613] = 8'b10000100;
DRAM[25614] = 8'b10000101;
DRAM[25615] = 8'b10000101;
DRAM[25616] = 8'b10000110;
DRAM[25617] = 8'b10000110;
DRAM[25618] = 8'b10000110;
DRAM[25619] = 8'b10000110;
DRAM[25620] = 8'b10000111;
DRAM[25621] = 8'b10001000;
DRAM[25622] = 8'b10001010;
DRAM[25623] = 8'b10001011;
DRAM[25624] = 8'b10001010;
DRAM[25625] = 8'b10001010;
DRAM[25626] = 8'b10011110;
DRAM[25627] = 8'b10100001;
DRAM[25628] = 8'b11001110;
DRAM[25629] = 8'b11000011;
DRAM[25630] = 8'b11011000;
DRAM[25631] = 8'b11100111;
DRAM[25632] = 8'b11010101;
DRAM[25633] = 8'b11000110;
DRAM[25634] = 8'b10110110;
DRAM[25635] = 8'b10111101;
DRAM[25636] = 8'b11000010;
DRAM[25637] = 8'b10100000;
DRAM[25638] = 8'b10010111;
DRAM[25639] = 8'b11001001;
DRAM[25640] = 8'b10100010;
DRAM[25641] = 8'b10101111;
DRAM[25642] = 8'b11001000;
DRAM[25643] = 8'b10101110;
DRAM[25644] = 8'b11000000;
DRAM[25645] = 8'b11001000;
DRAM[25646] = 8'b10110011;
DRAM[25647] = 8'b10110000;
DRAM[25648] = 8'b10111011;
DRAM[25649] = 8'b10101000;
DRAM[25650] = 8'b10110111;
DRAM[25651] = 8'b10111001;
DRAM[25652] = 8'b10110110;
DRAM[25653] = 8'b10101101;
DRAM[25654] = 8'b11001011;
DRAM[25655] = 8'b11001011;
DRAM[25656] = 8'b10111000;
DRAM[25657] = 8'b11001101;
DRAM[25658] = 8'b11010000;
DRAM[25659] = 8'b11000001;
DRAM[25660] = 8'b11100001;
DRAM[25661] = 8'b11100100;
DRAM[25662] = 8'b11100101;
DRAM[25663] = 8'b11100101;
DRAM[25664] = 8'b11011101;
DRAM[25665] = 8'b11011101;
DRAM[25666] = 8'b11011001;
DRAM[25667] = 8'b11001011;
DRAM[25668] = 8'b11100011;
DRAM[25669] = 8'b11100111;
DRAM[25670] = 8'b11001000;
DRAM[25671] = 8'b10111111;
DRAM[25672] = 8'b10110001;
DRAM[25673] = 8'b10110001;
DRAM[25674] = 8'b10110011;
DRAM[25675] = 8'b1110000;
DRAM[25676] = 8'b1100100;
DRAM[25677] = 8'b1101101;
DRAM[25678] = 8'b1101110;
DRAM[25679] = 8'b1101111;
DRAM[25680] = 8'b1111100;
DRAM[25681] = 8'b10001101;
DRAM[25682] = 8'b10011011;
DRAM[25683] = 8'b10100010;
DRAM[25684] = 8'b10101011;
DRAM[25685] = 8'b10111011;
DRAM[25686] = 8'b11000011;
DRAM[25687] = 8'b11000010;
DRAM[25688] = 8'b10111011;
DRAM[25689] = 8'b10110011;
DRAM[25690] = 8'b10110011;
DRAM[25691] = 8'b11000001;
DRAM[25692] = 8'b11001101;
DRAM[25693] = 8'b11010011;
DRAM[25694] = 8'b11011100;
DRAM[25695] = 8'b11100111;
DRAM[25696] = 8'b11100000;
DRAM[25697] = 8'b11011111;
DRAM[25698] = 8'b11011110;
DRAM[25699] = 8'b11011111;
DRAM[25700] = 8'b11011111;
DRAM[25701] = 8'b11011001;
DRAM[25702] = 8'b11001100;
DRAM[25703] = 8'b11000000;
DRAM[25704] = 8'b10111110;
DRAM[25705] = 8'b10111110;
DRAM[25706] = 8'b10110110;
DRAM[25707] = 8'b10110101;
DRAM[25708] = 8'b10111010;
DRAM[25709] = 8'b10110011;
DRAM[25710] = 8'b10101101;
DRAM[25711] = 8'b10110011;
DRAM[25712] = 8'b10101000;
DRAM[25713] = 8'b10111010;
DRAM[25714] = 8'b10101111;
DRAM[25715] = 8'b10001101;
DRAM[25716] = 8'b10110111;
DRAM[25717] = 8'b10010101;
DRAM[25718] = 8'b10010000;
DRAM[25719] = 8'b10101001;
DRAM[25720] = 8'b10100001;
DRAM[25721] = 8'b10101001;
DRAM[25722] = 8'b10100111;
DRAM[25723] = 8'b10011010;
DRAM[25724] = 8'b10010000;
DRAM[25725] = 8'b10011100;
DRAM[25726] = 8'b10101001;
DRAM[25727] = 8'b10011101;
DRAM[25728] = 8'b10001000;
DRAM[25729] = 8'b10010111;
DRAM[25730] = 8'b10011101;
DRAM[25731] = 8'b10010100;
DRAM[25732] = 8'b10001111;
DRAM[25733] = 8'b10011000;
DRAM[25734] = 8'b10100000;
DRAM[25735] = 8'b10100000;
DRAM[25736] = 8'b10100000;
DRAM[25737] = 8'b10100110;
DRAM[25738] = 8'b10101110;
DRAM[25739] = 8'b10110111;
DRAM[25740] = 8'b10101110;
DRAM[25741] = 8'b10100100;
DRAM[25742] = 8'b10011100;
DRAM[25743] = 8'b10011111;
DRAM[25744] = 8'b10100001;
DRAM[25745] = 8'b10011011;
DRAM[25746] = 8'b10010010;
DRAM[25747] = 8'b10010010;
DRAM[25748] = 8'b10100000;
DRAM[25749] = 8'b10011110;
DRAM[25750] = 8'b10001010;
DRAM[25751] = 8'b10000101;
DRAM[25752] = 8'b10001110;
DRAM[25753] = 8'b10001010;
DRAM[25754] = 8'b10000101;
DRAM[25755] = 8'b10000010;
DRAM[25756] = 8'b1111111;
DRAM[25757] = 8'b1111100;
DRAM[25758] = 8'b1110111;
DRAM[25759] = 8'b1110100;
DRAM[25760] = 8'b1101011;
DRAM[25761] = 8'b1100000;
DRAM[25762] = 8'b1100111;
DRAM[25763] = 8'b1110011;
DRAM[25764] = 8'b1101101;
DRAM[25765] = 8'b1010001;
DRAM[25766] = 8'b1001111;
DRAM[25767] = 8'b1011101;
DRAM[25768] = 8'b1011110;
DRAM[25769] = 8'b1100100;
DRAM[25770] = 8'b1110000;
DRAM[25771] = 8'b10000101;
DRAM[25772] = 8'b10010000;
DRAM[25773] = 8'b10001100;
DRAM[25774] = 8'b10010111;
DRAM[25775] = 8'b10110110;
DRAM[25776] = 8'b11000001;
DRAM[25777] = 8'b10111100;
DRAM[25778] = 8'b10111111;
DRAM[25779] = 8'b11000100;
DRAM[25780] = 8'b11000000;
DRAM[25781] = 8'b10111011;
DRAM[25782] = 8'b11001000;
DRAM[25783] = 8'b11011110;
DRAM[25784] = 8'b11100010;
DRAM[25785] = 8'b11101101;
DRAM[25786] = 8'b11101101;
DRAM[25787] = 8'b11101011;
DRAM[25788] = 8'b11101101;
DRAM[25789] = 8'b11100000;
DRAM[25790] = 8'b11001001;
DRAM[25791] = 8'b10111101;
DRAM[25792] = 8'b10101000;
DRAM[25793] = 8'b10100010;
DRAM[25794] = 8'b10001101;
DRAM[25795] = 8'b1111100;
DRAM[25796] = 8'b1100001;
DRAM[25797] = 8'b1101001;
DRAM[25798] = 8'b10010011;
DRAM[25799] = 8'b10001111;
DRAM[25800] = 8'b10011010;
DRAM[25801] = 8'b10101010;
DRAM[25802] = 8'b10110111;
DRAM[25803] = 8'b11010100;
DRAM[25804] = 8'b11110000;
DRAM[25805] = 8'b11101110;
DRAM[25806] = 8'b11100101;
DRAM[25807] = 8'b11100111;
DRAM[25808] = 8'b11101010;
DRAM[25809] = 8'b11011010;
DRAM[25810] = 8'b11100010;
DRAM[25811] = 8'b11001101;
DRAM[25812] = 8'b11001111;
DRAM[25813] = 8'b11011011;
DRAM[25814] = 8'b10111010;
DRAM[25815] = 8'b10100110;
DRAM[25816] = 8'b10101011;
DRAM[25817] = 8'b10110100;
DRAM[25818] = 8'b10011100;
DRAM[25819] = 8'b10100100;
DRAM[25820] = 8'b10100111;
DRAM[25821] = 8'b10010001;
DRAM[25822] = 8'b10011101;
DRAM[25823] = 8'b10100101;
DRAM[25824] = 8'b10011000;
DRAM[25825] = 8'b10011001;
DRAM[25826] = 8'b10010101;
DRAM[25827] = 8'b10011011;
DRAM[25828] = 8'b10101000;
DRAM[25829] = 8'b10111000;
DRAM[25830] = 8'b11001001;
DRAM[25831] = 8'b11001110;
DRAM[25832] = 8'b10101011;
DRAM[25833] = 8'b10010010;
DRAM[25834] = 8'b10010011;
DRAM[25835] = 8'b10010110;
DRAM[25836] = 8'b10000011;
DRAM[25837] = 8'b1110101;
DRAM[25838] = 8'b1110011;
DRAM[25839] = 8'b1110110;
DRAM[25840] = 8'b1101111;
DRAM[25841] = 8'b1101111;
DRAM[25842] = 8'b1101111;
DRAM[25843] = 8'b1101111;
DRAM[25844] = 8'b1101110;
DRAM[25845] = 8'b1101110;
DRAM[25846] = 8'b1101110;
DRAM[25847] = 8'b1101101;
DRAM[25848] = 8'b1101100;
DRAM[25849] = 8'b1101100;
DRAM[25850] = 8'b1101100;
DRAM[25851] = 8'b1101100;
DRAM[25852] = 8'b1101011;
DRAM[25853] = 8'b1101011;
DRAM[25854] = 8'b1101011;
DRAM[25855] = 8'b1101010;
DRAM[25856] = 8'b1111111;
DRAM[25857] = 8'b1111111;
DRAM[25858] = 8'b10000000;
DRAM[25859] = 8'b10000000;
DRAM[25860] = 8'b10000000;
DRAM[25861] = 8'b10000001;
DRAM[25862] = 8'b10000001;
DRAM[25863] = 8'b10000001;
DRAM[25864] = 8'b10000100;
DRAM[25865] = 8'b10000100;
DRAM[25866] = 8'b10000100;
DRAM[25867] = 8'b10000100;
DRAM[25868] = 8'b10000100;
DRAM[25869] = 8'b10000100;
DRAM[25870] = 8'b10000100;
DRAM[25871] = 8'b10000100;
DRAM[25872] = 8'b10000111;
DRAM[25873] = 8'b10000110;
DRAM[25874] = 8'b10000101;
DRAM[25875] = 8'b10000101;
DRAM[25876] = 8'b10000110;
DRAM[25877] = 8'b10001000;
DRAM[25878] = 8'b10001010;
DRAM[25879] = 8'b10001011;
DRAM[25880] = 8'b10000110;
DRAM[25881] = 8'b10010101;
DRAM[25882] = 8'b10010011;
DRAM[25883] = 8'b10010001;
DRAM[25884] = 8'b10111000;
DRAM[25885] = 8'b11001011;
DRAM[25886] = 8'b11010011;
DRAM[25887] = 8'b11011101;
DRAM[25888] = 8'b11010011;
DRAM[25889] = 8'b10111010;
DRAM[25890] = 8'b11000101;
DRAM[25891] = 8'b10111101;
DRAM[25892] = 8'b10100101;
DRAM[25893] = 8'b10101010;
DRAM[25894] = 8'b10101010;
DRAM[25895] = 8'b10100000;
DRAM[25896] = 8'b10101111;
DRAM[25897] = 8'b10110000;
DRAM[25898] = 8'b11000000;
DRAM[25899] = 8'b10110000;
DRAM[25900] = 8'b11000101;
DRAM[25901] = 8'b10101101;
DRAM[25902] = 8'b10101010;
DRAM[25903] = 8'b10111011;
DRAM[25904] = 8'b10111001;
DRAM[25905] = 8'b10100011;
DRAM[25906] = 8'b10111000;
DRAM[25907] = 8'b11000000;
DRAM[25908] = 8'b10101100;
DRAM[25909] = 8'b10100001;
DRAM[25910] = 8'b11001100;
DRAM[25911] = 8'b10111100;
DRAM[25912] = 8'b10111101;
DRAM[25913] = 8'b11001111;
DRAM[25914] = 8'b11001001;
DRAM[25915] = 8'b11000111;
DRAM[25916] = 8'b11010110;
DRAM[25917] = 8'b11100000;
DRAM[25918] = 8'b11011010;
DRAM[25919] = 8'b11100000;
DRAM[25920] = 8'b11011010;
DRAM[25921] = 8'b11010011;
DRAM[25922] = 8'b11010111;
DRAM[25923] = 8'b11000110;
DRAM[25924] = 8'b11011110;
DRAM[25925] = 8'b11100010;
DRAM[25926] = 8'b11001010;
DRAM[25927] = 8'b10110111;
DRAM[25928] = 8'b10100011;
DRAM[25929] = 8'b10100010;
DRAM[25930] = 8'b10011001;
DRAM[25931] = 8'b1011110;
DRAM[25932] = 8'b1011111;
DRAM[25933] = 8'b1101010;
DRAM[25934] = 8'b1110101;
DRAM[25935] = 8'b10000000;
DRAM[25936] = 8'b10000101;
DRAM[25937] = 8'b10010000;
DRAM[25938] = 8'b10011100;
DRAM[25939] = 8'b10100011;
DRAM[25940] = 8'b10101001;
DRAM[25941] = 8'b10110000;
DRAM[25942] = 8'b10110101;
DRAM[25943] = 8'b10110111;
DRAM[25944] = 8'b11000100;
DRAM[25945] = 8'b11000001;
DRAM[25946] = 8'b11000000;
DRAM[25947] = 8'b11000101;
DRAM[25948] = 8'b11001001;
DRAM[25949] = 8'b11001110;
DRAM[25950] = 8'b11010101;
DRAM[25951] = 8'b11011101;
DRAM[25952] = 8'b11011010;
DRAM[25953] = 8'b11011100;
DRAM[25954] = 8'b11011011;
DRAM[25955] = 8'b11011010;
DRAM[25956] = 8'b11011011;
DRAM[25957] = 8'b11011011;
DRAM[25958] = 8'b11010100;
DRAM[25959] = 8'b11001100;
DRAM[25960] = 8'b10110101;
DRAM[25961] = 8'b10110010;
DRAM[25962] = 8'b10100110;
DRAM[25963] = 8'b10100010;
DRAM[25964] = 8'b10100101;
DRAM[25965] = 8'b10100000;
DRAM[25966] = 8'b10011100;
DRAM[25967] = 8'b10100100;
DRAM[25968] = 8'b10011100;
DRAM[25969] = 8'b10010000;
DRAM[25970] = 8'b10101000;
DRAM[25971] = 8'b10001111;
DRAM[25972] = 8'b10011101;
DRAM[25973] = 8'b10000011;
DRAM[25974] = 8'b10011001;
DRAM[25975] = 8'b10001110;
DRAM[25976] = 8'b10011110;
DRAM[25977] = 8'b10110001;
DRAM[25978] = 8'b10100101;
DRAM[25979] = 8'b10011000;
DRAM[25980] = 8'b10011001;
DRAM[25981] = 8'b10100101;
DRAM[25982] = 8'b10110000;
DRAM[25983] = 8'b10011111;
DRAM[25984] = 8'b10001010;
DRAM[25985] = 8'b10011010;
DRAM[25986] = 8'b10011101;
DRAM[25987] = 8'b10010010;
DRAM[25988] = 8'b10010001;
DRAM[25989] = 8'b10011101;
DRAM[25990] = 8'b10011111;
DRAM[25991] = 8'b10010110;
DRAM[25992] = 8'b10100001;
DRAM[25993] = 8'b10100011;
DRAM[25994] = 8'b10100101;
DRAM[25995] = 8'b10110111;
DRAM[25996] = 8'b10101111;
DRAM[25997] = 8'b10101001;
DRAM[25998] = 8'b10011001;
DRAM[25999] = 8'b10011010;
DRAM[26000] = 8'b10010011;
DRAM[26001] = 8'b10011001;
DRAM[26002] = 8'b10100000;
DRAM[26003] = 8'b10010111;
DRAM[26004] = 8'b10011011;
DRAM[26005] = 8'b10011100;
DRAM[26006] = 8'b10001010;
DRAM[26007] = 8'b10001110;
DRAM[26008] = 8'b10010010;
DRAM[26009] = 8'b10001011;
DRAM[26010] = 8'b10001000;
DRAM[26011] = 8'b10001001;
DRAM[26012] = 8'b10000011;
DRAM[26013] = 8'b1110111;
DRAM[26014] = 8'b1110001;
DRAM[26015] = 8'b1110010;
DRAM[26016] = 8'b1101100;
DRAM[26017] = 8'b1011010;
DRAM[26018] = 8'b1011110;
DRAM[26019] = 8'b1100100;
DRAM[26020] = 8'b1101010;
DRAM[26021] = 8'b1010000;
DRAM[26022] = 8'b1010000;
DRAM[26023] = 8'b1010110;
DRAM[26024] = 8'b1100001;
DRAM[26025] = 8'b1110000;
DRAM[26026] = 8'b1110010;
DRAM[26027] = 8'b1101111;
DRAM[26028] = 8'b1110110;
DRAM[26029] = 8'b1111101;
DRAM[26030] = 8'b10000101;
DRAM[26031] = 8'b10010010;
DRAM[26032] = 8'b10001000;
DRAM[26033] = 8'b1111111;
DRAM[26034] = 8'b10001011;
DRAM[26035] = 8'b10100111;
DRAM[26036] = 8'b10110010;
DRAM[26037] = 8'b10101001;
DRAM[26038] = 8'b10101001;
DRAM[26039] = 8'b10110110;
DRAM[26040] = 8'b11010001;
DRAM[26041] = 8'b11011010;
DRAM[26042] = 8'b11011001;
DRAM[26043] = 8'b11010101;
DRAM[26044] = 8'b11011001;
DRAM[26045] = 8'b11010001;
DRAM[26046] = 8'b11000000;
DRAM[26047] = 8'b10111001;
DRAM[26048] = 8'b10100101;
DRAM[26049] = 8'b10011110;
DRAM[26050] = 8'b10000000;
DRAM[26051] = 8'b1110011;
DRAM[26052] = 8'b1010010;
DRAM[26053] = 8'b1010001;
DRAM[26054] = 8'b10000101;
DRAM[26055] = 8'b10001001;
DRAM[26056] = 8'b10010100;
DRAM[26057] = 8'b10101110;
DRAM[26058] = 8'b10110000;
DRAM[26059] = 8'b11001101;
DRAM[26060] = 8'b11110001;
DRAM[26061] = 8'b11101111;
DRAM[26062] = 8'b11101010;
DRAM[26063] = 8'b11101001;
DRAM[26064] = 8'b11100011;
DRAM[26065] = 8'b11011100;
DRAM[26066] = 8'b11010110;
DRAM[26067] = 8'b11011000;
DRAM[26068] = 8'b10111011;
DRAM[26069] = 8'b11011101;
DRAM[26070] = 8'b11000011;
DRAM[26071] = 8'b10100010;
DRAM[26072] = 8'b10101011;
DRAM[26073] = 8'b10110101;
DRAM[26074] = 8'b10100011;
DRAM[26075] = 8'b10100010;
DRAM[26076] = 8'b10101001;
DRAM[26077] = 8'b10010111;
DRAM[26078] = 8'b10010100;
DRAM[26079] = 8'b10100001;
DRAM[26080] = 8'b10010100;
DRAM[26081] = 8'b10011010;
DRAM[26082] = 8'b10010001;
DRAM[26083] = 8'b10011011;
DRAM[26084] = 8'b10101110;
DRAM[26085] = 8'b10111111;
DRAM[26086] = 8'b11001111;
DRAM[26087] = 8'b11000111;
DRAM[26088] = 8'b10110010;
DRAM[26089] = 8'b10000001;
DRAM[26090] = 8'b10000100;
DRAM[26091] = 8'b10010000;
DRAM[26092] = 8'b10000011;
DRAM[26093] = 8'b1110110;
DRAM[26094] = 8'b1101101;
DRAM[26095] = 8'b1110010;
DRAM[26096] = 8'b1110000;
DRAM[26097] = 8'b1110000;
DRAM[26098] = 8'b1110000;
DRAM[26099] = 8'b1101111;
DRAM[26100] = 8'b1101111;
DRAM[26101] = 8'b1101111;
DRAM[26102] = 8'b1101110;
DRAM[26103] = 8'b1101110;
DRAM[26104] = 8'b1101101;
DRAM[26105] = 8'b1101101;
DRAM[26106] = 8'b1101101;
DRAM[26107] = 8'b1101100;
DRAM[26108] = 8'b1101100;
DRAM[26109] = 8'b1101100;
DRAM[26110] = 8'b1101011;
DRAM[26111] = 8'b1101011;
DRAM[26112] = 8'b10000000;
DRAM[26113] = 8'b10000000;
DRAM[26114] = 8'b10000000;
DRAM[26115] = 8'b10000001;
DRAM[26116] = 8'b10000001;
DRAM[26117] = 8'b10000001;
DRAM[26118] = 8'b10000010;
DRAM[26119] = 8'b10000010;
DRAM[26120] = 8'b10000111;
DRAM[26121] = 8'b10000110;
DRAM[26122] = 8'b10000110;
DRAM[26123] = 8'b10000101;
DRAM[26124] = 8'b10000100;
DRAM[26125] = 8'b10000100;
DRAM[26126] = 8'b10000011;
DRAM[26127] = 8'b10000011;
DRAM[26128] = 8'b10000110;
DRAM[26129] = 8'b10000110;
DRAM[26130] = 8'b10000100;
DRAM[26131] = 8'b10000100;
DRAM[26132] = 8'b10000101;
DRAM[26133] = 8'b10000111;
DRAM[26134] = 8'b10001001;
DRAM[26135] = 8'b10001011;
DRAM[26136] = 8'b10001011;
DRAM[26137] = 8'b10011010;
DRAM[26138] = 8'b1111010;
DRAM[26139] = 8'b10010011;
DRAM[26140] = 8'b10101011;
DRAM[26141] = 8'b11010111;
DRAM[26142] = 8'b11000100;
DRAM[26143] = 8'b11010101;
DRAM[26144] = 8'b11010010;
DRAM[26145] = 8'b10111011;
DRAM[26146] = 8'b11000000;
DRAM[26147] = 8'b10100111;
DRAM[26148] = 8'b10011011;
DRAM[26149] = 8'b10111001;
DRAM[26150] = 8'b10101111;
DRAM[26151] = 8'b10001100;
DRAM[26152] = 8'b11000011;
DRAM[26153] = 8'b10101100;
DRAM[26154] = 8'b10101011;
DRAM[26155] = 8'b11000000;
DRAM[26156] = 8'b10110101;
DRAM[26157] = 8'b10011001;
DRAM[26158] = 8'b10101110;
DRAM[26159] = 8'b11000000;
DRAM[26160] = 8'b10100111;
DRAM[26161] = 8'b10101011;
DRAM[26162] = 8'b10110100;
DRAM[26163] = 8'b10101110;
DRAM[26164] = 8'b10101000;
DRAM[26165] = 8'b10100101;
DRAM[26166] = 8'b11001010;
DRAM[26167] = 8'b10110010;
DRAM[26168] = 8'b10111110;
DRAM[26169] = 8'b11001010;
DRAM[26170] = 8'b10111101;
DRAM[26171] = 8'b11001101;
DRAM[26172] = 8'b11001000;
DRAM[26173] = 8'b11011101;
DRAM[26174] = 8'b11010011;
DRAM[26175] = 8'b11100010;
DRAM[26176] = 8'b11011011;
DRAM[26177] = 8'b11001101;
DRAM[26178] = 8'b11011100;
DRAM[26179] = 8'b11001100;
DRAM[26180] = 8'b11011101;
DRAM[26181] = 8'b11100000;
DRAM[26182] = 8'b11001101;
DRAM[26183] = 8'b10101011;
DRAM[26184] = 8'b10101111;
DRAM[26185] = 8'b10100011;
DRAM[26186] = 8'b10000111;
DRAM[26187] = 8'b1010000;
DRAM[26188] = 8'b1011001;
DRAM[26189] = 8'b1011111;
DRAM[26190] = 8'b1101001;
DRAM[26191] = 8'b1110101;
DRAM[26192] = 8'b1111100;
DRAM[26193] = 8'b10000100;
DRAM[26194] = 8'b10010100;
DRAM[26195] = 8'b10100110;
DRAM[26196] = 8'b10110001;
DRAM[26197] = 8'b10110111;
DRAM[26198] = 8'b11000000;
DRAM[26199] = 8'b11001000;
DRAM[26200] = 8'b11001100;
DRAM[26201] = 8'b11010010;
DRAM[26202] = 8'b11010101;
DRAM[26203] = 8'b11010010;
DRAM[26204] = 8'b11001111;
DRAM[26205] = 8'b11010010;
DRAM[26206] = 8'b11010110;
DRAM[26207] = 8'b11010111;
DRAM[26208] = 8'b11100110;
DRAM[26209] = 8'b11100110;
DRAM[26210] = 8'b11100001;
DRAM[26211] = 8'b11011000;
DRAM[26212] = 8'b11010100;
DRAM[26213] = 8'b11010110;
DRAM[26214] = 8'b11010110;
DRAM[26215] = 8'b11010010;
DRAM[26216] = 8'b11000111;
DRAM[26217] = 8'b11000000;
DRAM[26218] = 8'b10101110;
DRAM[26219] = 8'b10100011;
DRAM[26220] = 8'b10100010;
DRAM[26221] = 8'b10011011;
DRAM[26222] = 8'b10011000;
DRAM[26223] = 8'b10100001;
DRAM[26224] = 8'b10100011;
DRAM[26225] = 8'b10010010;
DRAM[26226] = 8'b10011111;
DRAM[26227] = 8'b10010010;
DRAM[26228] = 8'b10010011;
DRAM[26229] = 8'b10001100;
DRAM[26230] = 8'b10011111;
DRAM[26231] = 8'b10010001;
DRAM[26232] = 8'b10001000;
DRAM[26233] = 8'b10100101;
DRAM[26234] = 8'b10010110;
DRAM[26235] = 8'b10010100;
DRAM[26236] = 8'b10011110;
DRAM[26237] = 8'b10011000;
DRAM[26238] = 8'b10011011;
DRAM[26239] = 8'b10010100;
DRAM[26240] = 8'b10010010;
DRAM[26241] = 8'b10010100;
DRAM[26242] = 8'b10010011;
DRAM[26243] = 8'b10010010;
DRAM[26244] = 8'b10010110;
DRAM[26245] = 8'b10011110;
DRAM[26246] = 8'b10011100;
DRAM[26247] = 8'b10010101;
DRAM[26248] = 8'b10100000;
DRAM[26249] = 8'b10011110;
DRAM[26250] = 8'b10011010;
DRAM[26251] = 8'b10110011;
DRAM[26252] = 8'b10101101;
DRAM[26253] = 8'b10101100;
DRAM[26254] = 8'b10010101;
DRAM[26255] = 8'b10010011;
DRAM[26256] = 8'b10010110;
DRAM[26257] = 8'b10010111;
DRAM[26258] = 8'b10100101;
DRAM[26259] = 8'b10011101;
DRAM[26260] = 8'b10011011;
DRAM[26261] = 8'b10010101;
DRAM[26262] = 8'b10000100;
DRAM[26263] = 8'b10011000;
DRAM[26264] = 8'b10000010;
DRAM[26265] = 8'b10000000;
DRAM[26266] = 8'b1111101;
DRAM[26267] = 8'b1111100;
DRAM[26268] = 8'b1111010;
DRAM[26269] = 8'b1110100;
DRAM[26270] = 8'b1101010;
DRAM[26271] = 8'b1100001;
DRAM[26272] = 8'b1101111;
DRAM[26273] = 8'b1011101;
DRAM[26274] = 8'b1100010;
DRAM[26275] = 8'b1011110;
DRAM[26276] = 8'b1100110;
DRAM[26277] = 8'b1001011;
DRAM[26278] = 8'b1001010;
DRAM[26279] = 8'b1001001;
DRAM[26280] = 8'b1010100;
DRAM[26281] = 8'b1010101;
DRAM[26282] = 8'b1001011;
DRAM[26283] = 8'b1001000;
DRAM[26284] = 8'b1010100;
DRAM[26285] = 8'b1011001;
DRAM[26286] = 8'b1010101;
DRAM[26287] = 8'b1010111;
DRAM[26288] = 8'b1111001;
DRAM[26289] = 8'b1110100;
DRAM[26290] = 8'b10000101;
DRAM[26291] = 8'b10101111;
DRAM[26292] = 8'b11001110;
DRAM[26293] = 8'b11001101;
DRAM[26294] = 8'b10111010;
DRAM[26295] = 8'b10101101;
DRAM[26296] = 8'b11001010;
DRAM[26297] = 8'b11010111;
DRAM[26298] = 8'b11010111;
DRAM[26299] = 8'b11010101;
DRAM[26300] = 8'b11011000;
DRAM[26301] = 8'b11010000;
DRAM[26302] = 8'b11000000;
DRAM[26303] = 8'b10111010;
DRAM[26304] = 8'b10101111;
DRAM[26305] = 8'b10101000;
DRAM[26306] = 8'b10001011;
DRAM[26307] = 8'b10000100;
DRAM[26308] = 8'b1011101;
DRAM[26309] = 8'b1001011;
DRAM[26310] = 8'b10000001;
DRAM[26311] = 8'b10001001;
DRAM[26312] = 8'b10010010;
DRAM[26313] = 8'b10110000;
DRAM[26314] = 8'b10101001;
DRAM[26315] = 8'b11000101;
DRAM[26316] = 8'b11110001;
DRAM[26317] = 8'b11110010;
DRAM[26318] = 8'b11101111;
DRAM[26319] = 8'b11101100;
DRAM[26320] = 8'b11100011;
DRAM[26321] = 8'b11011100;
DRAM[26322] = 8'b11010101;
DRAM[26323] = 8'b11101000;
DRAM[26324] = 8'b10110100;
DRAM[26325] = 8'b11001100;
DRAM[26326] = 8'b11001110;
DRAM[26327] = 8'b10101010;
DRAM[26328] = 8'b10100100;
DRAM[26329] = 8'b10101110;
DRAM[26330] = 8'b10101001;
DRAM[26331] = 8'b10011101;
DRAM[26332] = 8'b10101000;
DRAM[26333] = 8'b10011111;
DRAM[26334] = 8'b10001001;
DRAM[26335] = 8'b10011010;
DRAM[26336] = 8'b10010010;
DRAM[26337] = 8'b10011100;
DRAM[26338] = 8'b10010000;
DRAM[26339] = 8'b10011111;
DRAM[26340] = 8'b10110101;
DRAM[26341] = 8'b11000011;
DRAM[26342] = 8'b11001110;
DRAM[26343] = 8'b10111000;
DRAM[26344] = 8'b10110111;
DRAM[26345] = 8'b1111101;
DRAM[26346] = 8'b1111110;
DRAM[26347] = 8'b10000100;
DRAM[26348] = 8'b1110111;
DRAM[26349] = 8'b1110111;
DRAM[26350] = 8'b1101111;
DRAM[26351] = 8'b1110000;
DRAM[26352] = 8'b1110001;
DRAM[26353] = 8'b1110001;
DRAM[26354] = 8'b1110000;
DRAM[26355] = 8'b1110000;
DRAM[26356] = 8'b1110000;
DRAM[26357] = 8'b1101111;
DRAM[26358] = 8'b1101111;
DRAM[26359] = 8'b1101111;
DRAM[26360] = 8'b1101110;
DRAM[26361] = 8'b1101110;
DRAM[26362] = 8'b1101101;
DRAM[26363] = 8'b1101101;
DRAM[26364] = 8'b1101101;
DRAM[26365] = 8'b1101100;
DRAM[26366] = 8'b1101100;
DRAM[26367] = 8'b1101100;
DRAM[26368] = 8'b10000000;
DRAM[26369] = 8'b10000000;
DRAM[26370] = 8'b10000001;
DRAM[26371] = 8'b10000001;
DRAM[26372] = 8'b10000001;
DRAM[26373] = 8'b10000010;
DRAM[26374] = 8'b10000010;
DRAM[26375] = 8'b10000010;
DRAM[26376] = 8'b10001000;
DRAM[26377] = 8'b10001000;
DRAM[26378] = 8'b10000111;
DRAM[26379] = 8'b10000110;
DRAM[26380] = 8'b10000100;
DRAM[26381] = 8'b10000011;
DRAM[26382] = 8'b10000011;
DRAM[26383] = 8'b10000010;
DRAM[26384] = 8'b10000110;
DRAM[26385] = 8'b10000101;
DRAM[26386] = 8'b10000100;
DRAM[26387] = 8'b10000011;
DRAM[26388] = 8'b10000100;
DRAM[26389] = 8'b10000110;
DRAM[26390] = 8'b10001001;
DRAM[26391] = 8'b10001010;
DRAM[26392] = 8'b10001001;
DRAM[26393] = 8'b10001001;
DRAM[26394] = 8'b10001101;
DRAM[26395] = 8'b10010100;
DRAM[26396] = 8'b11000010;
DRAM[26397] = 8'b10110010;
DRAM[26398] = 8'b10111101;
DRAM[26399] = 8'b11100000;
DRAM[26400] = 8'b11011001;
DRAM[26401] = 8'b10111111;
DRAM[26402] = 8'b10110011;
DRAM[26403] = 8'b10101100;
DRAM[26404] = 8'b10110101;
DRAM[26405] = 8'b10100010;
DRAM[26406] = 8'b10001111;
DRAM[26407] = 8'b11000100;
DRAM[26408] = 8'b10100110;
DRAM[26409] = 8'b10101010;
DRAM[26410] = 8'b10101110;
DRAM[26411] = 8'b11001011;
DRAM[26412] = 8'b10011110;
DRAM[26413] = 8'b10100111;
DRAM[26414] = 8'b10111100;
DRAM[26415] = 8'b10011001;
DRAM[26416] = 8'b10011001;
DRAM[26417] = 8'b10111010;
DRAM[26418] = 8'b10110101;
DRAM[26419] = 8'b10011111;
DRAM[26420] = 8'b10101111;
DRAM[26421] = 8'b10110101;
DRAM[26422] = 8'b11010000;
DRAM[26423] = 8'b10110111;
DRAM[26424] = 8'b11000000;
DRAM[26425] = 8'b11001000;
DRAM[26426] = 8'b10110111;
DRAM[26427] = 8'b11010111;
DRAM[26428] = 8'b11000100;
DRAM[26429] = 8'b11100010;
DRAM[26430] = 8'b11011000;
DRAM[26431] = 8'b11101101;
DRAM[26432] = 8'b11011111;
DRAM[26433] = 8'b11001100;
DRAM[26434] = 8'b11100011;
DRAM[26435] = 8'b11010100;
DRAM[26436] = 8'b11100000;
DRAM[26437] = 8'b11100001;
DRAM[26438] = 8'b11010000;
DRAM[26439] = 8'b10100011;
DRAM[26440] = 8'b10100101;
DRAM[26441] = 8'b10010101;
DRAM[26442] = 8'b1110111;
DRAM[26443] = 8'b1001101;
DRAM[26444] = 8'b1100110;
DRAM[26445] = 8'b1101110;
DRAM[26446] = 8'b1111000;
DRAM[26447] = 8'b10000100;
DRAM[26448] = 8'b10010010;
DRAM[26449] = 8'b10010100;
DRAM[26450] = 8'b10011101;
DRAM[26451] = 8'b10101011;
DRAM[26452] = 8'b10101101;
DRAM[26453] = 8'b10100111;
DRAM[26454] = 8'b10101001;
DRAM[26455] = 8'b10110001;
DRAM[26456] = 8'b10100100;
DRAM[26457] = 8'b10110111;
DRAM[26458] = 8'b11000110;
DRAM[26459] = 8'b11001010;
DRAM[26460] = 8'b11001111;
DRAM[26461] = 8'b11011011;
DRAM[26462] = 8'b11100100;
DRAM[26463] = 8'b11100100;
DRAM[26464] = 8'b11011011;
DRAM[26465] = 8'b11100100;
DRAM[26466] = 8'b11100111;
DRAM[26467] = 8'b11100010;
DRAM[26468] = 8'b11011011;
DRAM[26469] = 8'b11010101;
DRAM[26470] = 8'b11001100;
DRAM[26471] = 8'b11000010;
DRAM[26472] = 8'b11000101;
DRAM[26473] = 8'b10111101;
DRAM[26474] = 8'b10101000;
DRAM[26475] = 8'b10011100;
DRAM[26476] = 8'b10011100;
DRAM[26477] = 8'b10010111;
DRAM[26478] = 8'b10010110;
DRAM[26479] = 8'b10100000;
DRAM[26480] = 8'b10100010;
DRAM[26481] = 8'b10100110;
DRAM[26482] = 8'b10000111;
DRAM[26483] = 8'b1110110;
DRAM[26484] = 8'b10000100;
DRAM[26485] = 8'b10000100;
DRAM[26486] = 8'b1111001;
DRAM[26487] = 8'b10001001;
DRAM[26488] = 8'b10000001;
DRAM[26489] = 8'b10100011;
DRAM[26490] = 8'b10010101;
DRAM[26491] = 8'b10100000;
DRAM[26492] = 8'b10101111;
DRAM[26493] = 8'b10010111;
DRAM[26494] = 8'b10010010;
DRAM[26495] = 8'b10011000;
DRAM[26496] = 8'b10011001;
DRAM[26497] = 8'b10001110;
DRAM[26498] = 8'b10001001;
DRAM[26499] = 8'b10010001;
DRAM[26500] = 8'b10011011;
DRAM[26501] = 8'b10011011;
DRAM[26502] = 8'b10011001;
DRAM[26503] = 8'b10011000;
DRAM[26504] = 8'b10100100;
DRAM[26505] = 8'b10011110;
DRAM[26506] = 8'b10010110;
DRAM[26507] = 8'b10110100;
DRAM[26508] = 8'b10110000;
DRAM[26509] = 8'b10110010;
DRAM[26510] = 8'b10010111;
DRAM[26511] = 8'b10010011;
DRAM[26512] = 8'b10100001;
DRAM[26513] = 8'b10010000;
DRAM[26514] = 8'b10011010;
DRAM[26515] = 8'b10011001;
DRAM[26516] = 8'b10011010;
DRAM[26517] = 8'b10001110;
DRAM[26518] = 8'b1111000;
DRAM[26519] = 8'b10010010;
DRAM[26520] = 8'b1111110;
DRAM[26521] = 8'b10000010;
DRAM[26522] = 8'b10000000;
DRAM[26523] = 8'b1111011;
DRAM[26524] = 8'b10000000;
DRAM[26525] = 8'b10000101;
DRAM[26526] = 8'b1111000;
DRAM[26527] = 8'b1100010;
DRAM[26528] = 8'b1101010;
DRAM[26529] = 8'b1100010;
DRAM[26530] = 8'b1101100;
DRAM[26531] = 8'b1011111;
DRAM[26532] = 8'b1011101;
DRAM[26533] = 8'b111100;
DRAM[26534] = 8'b111111;
DRAM[26535] = 8'b111111;
DRAM[26536] = 8'b1000000;
DRAM[26537] = 8'b1000110;
DRAM[26538] = 8'b1011000;
DRAM[26539] = 8'b1110011;
DRAM[26540] = 8'b1111100;
DRAM[26541] = 8'b1100111;
DRAM[26542] = 8'b1100010;
DRAM[26543] = 8'b1111001;
DRAM[26544] = 8'b10010000;
DRAM[26545] = 8'b10001110;
DRAM[26546] = 8'b10001111;
DRAM[26547] = 8'b10011000;
DRAM[26548] = 8'b10100101;
DRAM[26549] = 8'b10101111;
DRAM[26550] = 8'b10110001;
DRAM[26551] = 8'b10110000;
DRAM[26552] = 8'b10101001;
DRAM[26553] = 8'b10111101;
DRAM[26554] = 8'b11001010;
DRAM[26555] = 8'b11010010;
DRAM[26556] = 8'b11011100;
DRAM[26557] = 8'b11010111;
DRAM[26558] = 8'b11001000;
DRAM[26559] = 8'b11000010;
DRAM[26560] = 8'b10101100;
DRAM[26561] = 8'b10101000;
DRAM[26562] = 8'b10001110;
DRAM[26563] = 8'b10001100;
DRAM[26564] = 8'b1011100;
DRAM[26565] = 8'b111000;
DRAM[26566] = 8'b1100101;
DRAM[26567] = 8'b1101011;
DRAM[26568] = 8'b10010001;
DRAM[26569] = 8'b10110001;
DRAM[26570] = 8'b10100101;
DRAM[26571] = 8'b11000001;
DRAM[26572] = 8'b11110001;
DRAM[26573] = 8'b11110100;
DRAM[26574] = 8'b11110011;
DRAM[26575] = 8'b11101111;
DRAM[26576] = 8'b11101000;
DRAM[26577] = 8'b11011011;
DRAM[26578] = 8'b11011011;
DRAM[26579] = 8'b11110110;
DRAM[26580] = 8'b10110110;
DRAM[26581] = 8'b10111011;
DRAM[26582] = 8'b11010111;
DRAM[26583] = 8'b10110101;
DRAM[26584] = 8'b10011011;
DRAM[26585] = 8'b10100101;
DRAM[26586] = 8'b10101010;
DRAM[26587] = 8'b10010111;
DRAM[26588] = 8'b10100100;
DRAM[26589] = 8'b10100011;
DRAM[26590] = 8'b10000000;
DRAM[26591] = 8'b10010101;
DRAM[26592] = 8'b10010011;
DRAM[26593] = 8'b10011111;
DRAM[26594] = 8'b10010010;
DRAM[26595] = 8'b10100011;
DRAM[26596] = 8'b10111010;
DRAM[26597] = 8'b11000100;
DRAM[26598] = 8'b11001001;
DRAM[26599] = 8'b10101010;
DRAM[26600] = 8'b10110110;
DRAM[26601] = 8'b1111101;
DRAM[26602] = 8'b1111101;
DRAM[26603] = 8'b1111001;
DRAM[26604] = 8'b1101100;
DRAM[26605] = 8'b1111001;
DRAM[26606] = 8'b1110101;
DRAM[26607] = 8'b1110001;
DRAM[26608] = 8'b1110001;
DRAM[26609] = 8'b1110001;
DRAM[26610] = 8'b1110001;
DRAM[26611] = 8'b1110000;
DRAM[26612] = 8'b1110000;
DRAM[26613] = 8'b1110000;
DRAM[26614] = 8'b1101111;
DRAM[26615] = 8'b1101111;
DRAM[26616] = 8'b1101110;
DRAM[26617] = 8'b1101110;
DRAM[26618] = 8'b1101110;
DRAM[26619] = 8'b1101101;
DRAM[26620] = 8'b1101101;
DRAM[26621] = 8'b1101101;
DRAM[26622] = 8'b1101100;
DRAM[26623] = 8'b1101100;
DRAM[26624] = 8'b10000011;
DRAM[26625] = 8'b10000011;
DRAM[26626] = 8'b10000100;
DRAM[26627] = 8'b10000100;
DRAM[26628] = 8'b10000100;
DRAM[26629] = 8'b10000101;
DRAM[26630] = 8'b10000101;
DRAM[26631] = 8'b10000101;
DRAM[26632] = 8'b10000100;
DRAM[26633] = 8'b10000100;
DRAM[26634] = 8'b10000100;
DRAM[26635] = 8'b10000100;
DRAM[26636] = 8'b10000100;
DRAM[26637] = 8'b10000100;
DRAM[26638] = 8'b10000011;
DRAM[26639] = 8'b10000011;
DRAM[26640] = 8'b10000110;
DRAM[26641] = 8'b10000110;
DRAM[26642] = 8'b10000110;
DRAM[26643] = 8'b10000111;
DRAM[26644] = 8'b10000111;
DRAM[26645] = 8'b10000111;
DRAM[26646] = 8'b10001000;
DRAM[26647] = 8'b10001000;
DRAM[26648] = 8'b10010000;
DRAM[26649] = 8'b10000101;
DRAM[26650] = 8'b10000110;
DRAM[26651] = 8'b10011001;
DRAM[26652] = 8'b10101001;
DRAM[26653] = 8'b10110000;
DRAM[26654] = 8'b10111100;
DRAM[26655] = 8'b11001011;
DRAM[26656] = 8'b11010011;
DRAM[26657] = 8'b11001100;
DRAM[26658] = 8'b10110111;
DRAM[26659] = 8'b11000001;
DRAM[26660] = 8'b10110011;
DRAM[26661] = 8'b10010110;
DRAM[26662] = 8'b10101100;
DRAM[26663] = 8'b10111100;
DRAM[26664] = 8'b10100000;
DRAM[26665] = 8'b10100011;
DRAM[26666] = 8'b10111010;
DRAM[26667] = 8'b10010110;
DRAM[26668] = 8'b10100111;
DRAM[26669] = 8'b10110110;
DRAM[26670] = 8'b10101001;
DRAM[26671] = 8'b10010010;
DRAM[26672] = 8'b10110111;
DRAM[26673] = 8'b11000000;
DRAM[26674] = 8'b10100111;
DRAM[26675] = 8'b10110001;
DRAM[26676] = 8'b10110111;
DRAM[26677] = 8'b10111100;
DRAM[26678] = 8'b10110001;
DRAM[26679] = 8'b11010100;
DRAM[26680] = 8'b10101111;
DRAM[26681] = 8'b10111001;
DRAM[26682] = 8'b11001110;
DRAM[26683] = 8'b11001000;
DRAM[26684] = 8'b11001100;
DRAM[26685] = 8'b11110111;
DRAM[26686] = 8'b11010011;
DRAM[26687] = 8'b11100010;
DRAM[26688] = 8'b11011100;
DRAM[26689] = 8'b11011011;
DRAM[26690] = 8'b11101001;
DRAM[26691] = 8'b11001011;
DRAM[26692] = 8'b11100111;
DRAM[26693] = 8'b11011110;
DRAM[26694] = 8'b10111101;
DRAM[26695] = 8'b10110101;
DRAM[26696] = 8'b10010110;
DRAM[26697] = 8'b10010111;
DRAM[26698] = 8'b1110100;
DRAM[26699] = 8'b1000000;
DRAM[26700] = 8'b1011011;
DRAM[26701] = 8'b1100000;
DRAM[26702] = 8'b1101111;
DRAM[26703] = 8'b1111100;
DRAM[26704] = 8'b10001100;
DRAM[26705] = 8'b10011010;
DRAM[26706] = 8'b10100011;
DRAM[26707] = 8'b10101011;
DRAM[26708] = 8'b10110111;
DRAM[26709] = 8'b10111001;
DRAM[26710] = 8'b10111001;
DRAM[26711] = 8'b11000010;
DRAM[26712] = 8'b11000011;
DRAM[26713] = 8'b11001100;
DRAM[26714] = 8'b11010111;
DRAM[26715] = 8'b11011110;
DRAM[26716] = 8'b11100010;
DRAM[26717] = 8'b11100111;
DRAM[26718] = 8'b11101100;
DRAM[26719] = 8'b11110000;
DRAM[26720] = 8'b11100011;
DRAM[26721] = 8'b11100000;
DRAM[26722] = 8'b11011100;
DRAM[26723] = 8'b11011011;
DRAM[26724] = 8'b11011100;
DRAM[26725] = 8'b11011011;
DRAM[26726] = 8'b11010011;
DRAM[26727] = 8'b11001010;
DRAM[26728] = 8'b10110011;
DRAM[26729] = 8'b10101100;
DRAM[26730] = 8'b10111100;
DRAM[26731] = 8'b10101010;
DRAM[26732] = 8'b10011100;
DRAM[26733] = 8'b10010110;
DRAM[26734] = 8'b1110110;
DRAM[26735] = 8'b1110100;
DRAM[26736] = 8'b10011011;
DRAM[26737] = 8'b10010110;
DRAM[26738] = 8'b10001010;
DRAM[26739] = 8'b10000010;
DRAM[26740] = 8'b10000000;
DRAM[26741] = 8'b1111011;
DRAM[26742] = 8'b1111111;
DRAM[26743] = 8'b10001111;
DRAM[26744] = 8'b1111111;
DRAM[26745] = 8'b10010111;
DRAM[26746] = 8'b10011011;
DRAM[26747] = 8'b10001011;
DRAM[26748] = 8'b10100110;
DRAM[26749] = 8'b10010111;
DRAM[26750] = 8'b10001111;
DRAM[26751] = 8'b10010110;
DRAM[26752] = 8'b10011110;
DRAM[26753] = 8'b1111001;
DRAM[26754] = 8'b10011101;
DRAM[26755] = 8'b10011011;
DRAM[26756] = 8'b10000101;
DRAM[26757] = 8'b10010100;
DRAM[26758] = 8'b10010011;
DRAM[26759] = 8'b10100110;
DRAM[26760] = 8'b10100101;
DRAM[26761] = 8'b10011101;
DRAM[26762] = 8'b10100001;
DRAM[26763] = 8'b10100011;
DRAM[26764] = 8'b10100100;
DRAM[26765] = 8'b10110101;
DRAM[26766] = 8'b10110001;
DRAM[26767] = 8'b10001110;
DRAM[26768] = 8'b10111011;
DRAM[26769] = 8'b10010100;
DRAM[26770] = 8'b10100010;
DRAM[26771] = 8'b10100001;
DRAM[26772] = 8'b10010101;
DRAM[26773] = 8'b1111101;
DRAM[26774] = 8'b10010011;
DRAM[26775] = 8'b10001110;
DRAM[26776] = 8'b10010110;
DRAM[26777] = 8'b1111000;
DRAM[26778] = 8'b1110110;
DRAM[26779] = 8'b10000011;
DRAM[26780] = 8'b1111101;
DRAM[26781] = 8'b1110111;
DRAM[26782] = 8'b1110011;
DRAM[26783] = 8'b1100110;
DRAM[26784] = 8'b1101000;
DRAM[26785] = 8'b1100001;
DRAM[26786] = 8'b1100001;
DRAM[26787] = 8'b1100111;
DRAM[26788] = 8'b1011111;
DRAM[26789] = 8'b1000110;
DRAM[26790] = 8'b101101;
DRAM[26791] = 8'b100001;
DRAM[26792] = 8'b1000001;
DRAM[26793] = 8'b1000100;
DRAM[26794] = 8'b1001110;
DRAM[26795] = 8'b1111011;
DRAM[26796] = 8'b1011011;
DRAM[26797] = 8'b10100111;
DRAM[26798] = 8'b11010010;
DRAM[26799] = 8'b10101010;
DRAM[26800] = 8'b10101010;
DRAM[26801] = 8'b10011111;
DRAM[26802] = 8'b10000111;
DRAM[26803] = 8'b10100110;
DRAM[26804] = 8'b10111001;
DRAM[26805] = 8'b10100011;
DRAM[26806] = 8'b10100111;
DRAM[26807] = 8'b10101001;
DRAM[26808] = 8'b10101011;
DRAM[26809] = 8'b10111111;
DRAM[26810] = 8'b11000101;
DRAM[26811] = 8'b10111011;
DRAM[26812] = 8'b10111111;
DRAM[26813] = 8'b11001101;
DRAM[26814] = 8'b11000101;
DRAM[26815] = 8'b10101100;
DRAM[26816] = 8'b10010111;
DRAM[26817] = 8'b10010110;
DRAM[26818] = 8'b10000101;
DRAM[26819] = 8'b1101001;
DRAM[26820] = 8'b1100001;
DRAM[26821] = 8'b1001110;
DRAM[26822] = 8'b1000110;
DRAM[26823] = 8'b1110111;
DRAM[26824] = 8'b10001101;
DRAM[26825] = 8'b10011011;
DRAM[26826] = 8'b10100001;
DRAM[26827] = 8'b11000011;
DRAM[26828] = 8'b11101001;
DRAM[26829] = 8'b11110100;
DRAM[26830] = 8'b11111001;
DRAM[26831] = 8'b11110111;
DRAM[26832] = 8'b11101011;
DRAM[26833] = 8'b11101001;
DRAM[26834] = 8'b11101111;
DRAM[26835] = 8'b11011011;
DRAM[26836] = 8'b11100101;
DRAM[26837] = 8'b10111010;
DRAM[26838] = 8'b11010001;
DRAM[26839] = 8'b10101010;
DRAM[26840] = 8'b10100011;
DRAM[26841] = 8'b10101000;
DRAM[26842] = 8'b10100100;
DRAM[26843] = 8'b10011110;
DRAM[26844] = 8'b10001101;
DRAM[26845] = 8'b10100000;
DRAM[26846] = 8'b10001000;
DRAM[26847] = 8'b10000101;
DRAM[26848] = 8'b10010111;
DRAM[26849] = 8'b10011010;
DRAM[26850] = 8'b10011110;
DRAM[26851] = 8'b10101011;
DRAM[26852] = 8'b11000100;
DRAM[26853] = 8'b11000101;
DRAM[26854] = 8'b10100110;
DRAM[26855] = 8'b10101000;
DRAM[26856] = 8'b10010101;
DRAM[26857] = 8'b10000110;
DRAM[26858] = 8'b1111000;
DRAM[26859] = 8'b1110101;
DRAM[26860] = 8'b1110111;
DRAM[26861] = 8'b1110111;
DRAM[26862] = 8'b1110110;
DRAM[26863] = 8'b1110111;
DRAM[26864] = 8'b1110011;
DRAM[26865] = 8'b1110010;
DRAM[26866] = 8'b1110000;
DRAM[26867] = 8'b1110000;
DRAM[26868] = 8'b1110010;
DRAM[26869] = 8'b1110010;
DRAM[26870] = 8'b1110000;
DRAM[26871] = 8'b1101111;
DRAM[26872] = 8'b1110000;
DRAM[26873] = 8'b1110000;
DRAM[26874] = 8'b1101111;
DRAM[26875] = 8'b1101110;
DRAM[26876] = 8'b1101110;
DRAM[26877] = 8'b1101101;
DRAM[26878] = 8'b1101100;
DRAM[26879] = 8'b1101100;
DRAM[26880] = 8'b10000001;
DRAM[26881] = 8'b10000010;
DRAM[26882] = 8'b10000010;
DRAM[26883] = 8'b10000010;
DRAM[26884] = 8'b10000011;
DRAM[26885] = 8'b10000011;
DRAM[26886] = 8'b10000011;
DRAM[26887] = 8'b10000100;
DRAM[26888] = 8'b10000101;
DRAM[26889] = 8'b10000101;
DRAM[26890] = 8'b10000101;
DRAM[26891] = 8'b10000101;
DRAM[26892] = 8'b10000101;
DRAM[26893] = 8'b10000101;
DRAM[26894] = 8'b10000101;
DRAM[26895] = 8'b10000100;
DRAM[26896] = 8'b10000111;
DRAM[26897] = 8'b10000111;
DRAM[26898] = 8'b10000111;
DRAM[26899] = 8'b10000111;
DRAM[26900] = 8'b10001000;
DRAM[26901] = 8'b10001000;
DRAM[26902] = 8'b10001001;
DRAM[26903] = 8'b10001001;
DRAM[26904] = 8'b10001100;
DRAM[26905] = 8'b10001011;
DRAM[26906] = 8'b10010000;
DRAM[26907] = 8'b10011100;
DRAM[26908] = 8'b10100011;
DRAM[26909] = 8'b10101001;
DRAM[26910] = 8'b10110110;
DRAM[26911] = 8'b11000101;
DRAM[26912] = 8'b11001000;
DRAM[26913] = 8'b11010101;
DRAM[26914] = 8'b11000010;
DRAM[26915] = 8'b10110111;
DRAM[26916] = 8'b10101001;
DRAM[26917] = 8'b10100010;
DRAM[26918] = 8'b10110000;
DRAM[26919] = 8'b10100110;
DRAM[26920] = 8'b10100110;
DRAM[26921] = 8'b10011110;
DRAM[26922] = 8'b10100111;
DRAM[26923] = 8'b10100100;
DRAM[26924] = 8'b10100101;
DRAM[26925] = 8'b10101111;
DRAM[26926] = 8'b10011010;
DRAM[26927] = 8'b10011011;
DRAM[26928] = 8'b10111010;
DRAM[26929] = 8'b10111001;
DRAM[26930] = 8'b10100110;
DRAM[26931] = 8'b10101001;
DRAM[26932] = 8'b10101111;
DRAM[26933] = 8'b10110000;
DRAM[26934] = 8'b10101101;
DRAM[26935] = 8'b11000110;
DRAM[26936] = 8'b10111011;
DRAM[26937] = 8'b11000001;
DRAM[26938] = 8'b11010010;
DRAM[26939] = 8'b11001111;
DRAM[26940] = 8'b11010111;
DRAM[26941] = 8'b11110000;
DRAM[26942] = 8'b11011011;
DRAM[26943] = 8'b11100100;
DRAM[26944] = 8'b11110001;
DRAM[26945] = 8'b11011000;
DRAM[26946] = 8'b11011100;
DRAM[26947] = 8'b11010001;
DRAM[26948] = 8'b11101010;
DRAM[26949] = 8'b11010010;
DRAM[26950] = 8'b10110011;
DRAM[26951] = 8'b10111000;
DRAM[26952] = 8'b10011001;
DRAM[26953] = 8'b10010011;
DRAM[26954] = 8'b1101110;
DRAM[26955] = 8'b1001100;
DRAM[26956] = 8'b1100100;
DRAM[26957] = 8'b1101011;
DRAM[26958] = 8'b1110001;
DRAM[26959] = 8'b1111111;
DRAM[26960] = 8'b10000011;
DRAM[26961] = 8'b10011001;
DRAM[26962] = 8'b10100110;
DRAM[26963] = 8'b10100111;
DRAM[26964] = 8'b10101010;
DRAM[26965] = 8'b10101111;
DRAM[26966] = 8'b11000000;
DRAM[26967] = 8'b11011001;
DRAM[26968] = 8'b11011001;
DRAM[26969] = 8'b11010010;
DRAM[26970] = 8'b11010100;
DRAM[26971] = 8'b11100000;
DRAM[26972] = 8'b11101011;
DRAM[26973] = 8'b11101011;
DRAM[26974] = 8'b11101000;
DRAM[26975] = 8'b11101000;
DRAM[26976] = 8'b11100100;
DRAM[26977] = 8'b11101101;
DRAM[26978] = 8'b11101010;
DRAM[26979] = 8'b11010100;
DRAM[26980] = 8'b11000001;
DRAM[26981] = 8'b10111011;
DRAM[26982] = 8'b10111000;
DRAM[26983] = 8'b10110010;
DRAM[26984] = 8'b10110010;
DRAM[26985] = 8'b10100111;
DRAM[26986] = 8'b10100100;
DRAM[26987] = 8'b10010101;
DRAM[26988] = 8'b10001011;
DRAM[26989] = 8'b10001001;
DRAM[26990] = 8'b10000001;
DRAM[26991] = 8'b10000111;
DRAM[26992] = 8'b1110000;
DRAM[26993] = 8'b10000010;
DRAM[26994] = 8'b10001101;
DRAM[26995] = 8'b10000001;
DRAM[26996] = 8'b1101100;
DRAM[26997] = 8'b1100110;
DRAM[26998] = 8'b1110000;
DRAM[26999] = 8'b1111010;
DRAM[27000] = 8'b1111000;
DRAM[27001] = 8'b10001111;
DRAM[27002] = 8'b10010110;
DRAM[27003] = 8'b10000101;
DRAM[27004] = 8'b10011100;
DRAM[27005] = 8'b10001110;
DRAM[27006] = 8'b10001101;
DRAM[27007] = 8'b10011000;
DRAM[27008] = 8'b10010100;
DRAM[27009] = 8'b10000011;
DRAM[27010] = 8'b10100011;
DRAM[27011] = 8'b10010110;
DRAM[27012] = 8'b10001001;
DRAM[27013] = 8'b10011111;
DRAM[27014] = 8'b10011000;
DRAM[27015] = 8'b10011110;
DRAM[27016] = 8'b10011011;
DRAM[27017] = 8'b10011111;
DRAM[27018] = 8'b10100110;
DRAM[27019] = 8'b10101000;
DRAM[27020] = 8'b10101101;
DRAM[27021] = 8'b10110111;
DRAM[27022] = 8'b10101110;
DRAM[27023] = 8'b10010011;
DRAM[27024] = 8'b10110110;
DRAM[27025] = 8'b10100010;
DRAM[27026] = 8'b10100011;
DRAM[27027] = 8'b10101100;
DRAM[27028] = 8'b10010100;
DRAM[27029] = 8'b10001000;
DRAM[27030] = 8'b10001000;
DRAM[27031] = 8'b10000111;
DRAM[27032] = 8'b10011110;
DRAM[27033] = 8'b10001000;
DRAM[27034] = 8'b10000001;
DRAM[27035] = 8'b10000111;
DRAM[27036] = 8'b10000100;
DRAM[27037] = 8'b1111010;
DRAM[27038] = 8'b1110010;
DRAM[27039] = 8'b1101010;
DRAM[27040] = 8'b1101001;
DRAM[27041] = 8'b1011101;
DRAM[27042] = 8'b1011001;
DRAM[27043] = 8'b1011101;
DRAM[27044] = 8'b1010010;
DRAM[27045] = 8'b110101;
DRAM[27046] = 8'b11111;
DRAM[27047] = 8'b11010;
DRAM[27048] = 8'b101100;
DRAM[27049] = 8'b11010;
DRAM[27050] = 8'b10110;
DRAM[27051] = 8'b1000101;
DRAM[27052] = 8'b1101001;
DRAM[27053] = 8'b1100110;
DRAM[27054] = 8'b1101001;
DRAM[27055] = 8'b10111000;
DRAM[27056] = 8'b10101010;
DRAM[27057] = 8'b10110001;
DRAM[27058] = 8'b10101010;
DRAM[27059] = 8'b10111010;
DRAM[27060] = 8'b11000000;
DRAM[27061] = 8'b10110101;
DRAM[27062] = 8'b10110101;
DRAM[27063] = 8'b10100000;
DRAM[27064] = 8'b10011001;
DRAM[27065] = 8'b10101000;
DRAM[27066] = 8'b10111111;
DRAM[27067] = 8'b11001011;
DRAM[27068] = 8'b10111100;
DRAM[27069] = 8'b10100110;
DRAM[27070] = 8'b10100110;
DRAM[27071] = 8'b10110101;
DRAM[27072] = 8'b10011001;
DRAM[27073] = 8'b10010111;
DRAM[27074] = 8'b10001011;
DRAM[27075] = 8'b1110011;
DRAM[27076] = 8'b1101011;
DRAM[27077] = 8'b1010110;
DRAM[27078] = 8'b1001000;
DRAM[27079] = 8'b1110000;
DRAM[27080] = 8'b10000111;
DRAM[27081] = 8'b10011001;
DRAM[27082] = 8'b10101101;
DRAM[27083] = 8'b10101000;
DRAM[27084] = 8'b11001101;
DRAM[27085] = 8'b11111101;
DRAM[27086] = 8'b11110110;
DRAM[27087] = 8'b11110010;
DRAM[27088] = 8'b11111001;
DRAM[27089] = 8'b11101001;
DRAM[27090] = 8'b11101100;
DRAM[27091] = 8'b11011110;
DRAM[27092] = 8'b11011101;
DRAM[27093] = 8'b10111100;
DRAM[27094] = 8'b11001011;
DRAM[27095] = 8'b10111110;
DRAM[27096] = 8'b10101100;
DRAM[27097] = 8'b10011100;
DRAM[27098] = 8'b10100001;
DRAM[27099] = 8'b10011011;
DRAM[27100] = 8'b10011100;
DRAM[27101] = 8'b10010110;
DRAM[27102] = 8'b10001001;
DRAM[27103] = 8'b10001101;
DRAM[27104] = 8'b10010100;
DRAM[27105] = 8'b10011010;
DRAM[27106] = 8'b10011110;
DRAM[27107] = 8'b10110100;
DRAM[27108] = 8'b11000110;
DRAM[27109] = 8'b10111011;
DRAM[27110] = 8'b10101000;
DRAM[27111] = 8'b10100010;
DRAM[27112] = 8'b10001011;
DRAM[27113] = 8'b1111110;
DRAM[27114] = 8'b1110011;
DRAM[27115] = 8'b1110010;
DRAM[27116] = 8'b1110110;
DRAM[27117] = 8'b1110111;
DRAM[27118] = 8'b1110111;
DRAM[27119] = 8'b1111000;
DRAM[27120] = 8'b1110011;
DRAM[27121] = 8'b1110010;
DRAM[27122] = 8'b1110000;
DRAM[27123] = 8'b1110001;
DRAM[27124] = 8'b1110010;
DRAM[27125] = 8'b1110010;
DRAM[27126] = 8'b1110001;
DRAM[27127] = 8'b1101111;
DRAM[27128] = 8'b1110000;
DRAM[27129] = 8'b1110000;
DRAM[27130] = 8'b1101111;
DRAM[27131] = 8'b1101111;
DRAM[27132] = 8'b1101110;
DRAM[27133] = 8'b1101101;
DRAM[27134] = 8'b1101100;
DRAM[27135] = 8'b1101100;
DRAM[27136] = 8'b10000000;
DRAM[27137] = 8'b10000000;
DRAM[27138] = 8'b10000001;
DRAM[27139] = 8'b10000001;
DRAM[27140] = 8'b10000001;
DRAM[27141] = 8'b10000010;
DRAM[27142] = 8'b10000010;
DRAM[27143] = 8'b10000010;
DRAM[27144] = 8'b10000110;
DRAM[27145] = 8'b10000110;
DRAM[27146] = 8'b10000110;
DRAM[27147] = 8'b10000110;
DRAM[27148] = 8'b10000110;
DRAM[27149] = 8'b10000110;
DRAM[27150] = 8'b10000110;
DRAM[27151] = 8'b10000110;
DRAM[27152] = 8'b10001000;
DRAM[27153] = 8'b10001000;
DRAM[27154] = 8'b10001000;
DRAM[27155] = 8'b10001001;
DRAM[27156] = 8'b10001001;
DRAM[27157] = 8'b10001001;
DRAM[27158] = 8'b10001010;
DRAM[27159] = 8'b10001010;
DRAM[27160] = 8'b10001000;
DRAM[27161] = 8'b10010000;
DRAM[27162] = 8'b10011001;
DRAM[27163] = 8'b10011010;
DRAM[27164] = 8'b10011001;
DRAM[27165] = 8'b10011111;
DRAM[27166] = 8'b10101110;
DRAM[27167] = 8'b10111011;
DRAM[27168] = 8'b10111000;
DRAM[27169] = 8'b11011000;
DRAM[27170] = 8'b11001101;
DRAM[27171] = 8'b10110000;
DRAM[27172] = 8'b10100100;
DRAM[27173] = 8'b10110001;
DRAM[27174] = 8'b10110101;
DRAM[27175] = 8'b10010101;
DRAM[27176] = 8'b10101011;
DRAM[27177] = 8'b10011001;
DRAM[27178] = 8'b10010110;
DRAM[27179] = 8'b10110010;
DRAM[27180] = 8'b10100011;
DRAM[27181] = 8'b10100011;
DRAM[27182] = 8'b10001110;
DRAM[27183] = 8'b10101000;
DRAM[27184] = 8'b10111001;
DRAM[27185] = 8'b10101100;
DRAM[27186] = 8'b10100110;
DRAM[27187] = 8'b10100010;
DRAM[27188] = 8'b10101010;
DRAM[27189] = 8'b10100111;
DRAM[27190] = 8'b10110001;
DRAM[27191] = 8'b10111011;
DRAM[27192] = 8'b11000010;
DRAM[27193] = 8'b11000010;
DRAM[27194] = 8'b11001101;
DRAM[27195] = 8'b11001111;
DRAM[27196] = 8'b11011100;
DRAM[27197] = 8'b11011101;
DRAM[27198] = 8'b11011110;
DRAM[27199] = 8'b11011101;
DRAM[27200] = 8'b11101110;
DRAM[27201] = 8'b11010101;
DRAM[27202] = 8'b11010101;
DRAM[27203] = 8'b11010110;
DRAM[27204] = 8'b11101001;
DRAM[27205] = 8'b11010000;
DRAM[27206] = 8'b10101110;
DRAM[27207] = 8'b10101010;
DRAM[27208] = 8'b10100010;
DRAM[27209] = 8'b10001011;
DRAM[27210] = 8'b1011001;
DRAM[27211] = 8'b1001101;
DRAM[27212] = 8'b1011101;
DRAM[27213] = 8'b1101011;
DRAM[27214] = 8'b1101001;
DRAM[27215] = 8'b1111110;
DRAM[27216] = 8'b10001101;
DRAM[27217] = 8'b10011100;
DRAM[27218] = 8'b10100111;
DRAM[27219] = 8'b10110100;
DRAM[27220] = 8'b11000011;
DRAM[27221] = 8'b11000111;
DRAM[27222] = 8'b11000111;
DRAM[27223] = 8'b11001110;
DRAM[27224] = 8'b11001111;
DRAM[27225] = 8'b11000111;
DRAM[27226] = 8'b11000111;
DRAM[27227] = 8'b11010011;
DRAM[27228] = 8'b11011011;
DRAM[27229] = 8'b11011000;
DRAM[27230] = 8'b11010110;
DRAM[27231] = 8'b11011001;
DRAM[27232] = 8'b11100100;
DRAM[27233] = 8'b11100111;
DRAM[27234] = 8'b11011111;
DRAM[27235] = 8'b11010000;
DRAM[27236] = 8'b11001001;
DRAM[27237] = 8'b11000101;
DRAM[27238] = 8'b10110010;
DRAM[27239] = 8'b10011010;
DRAM[27240] = 8'b10100101;
DRAM[27241] = 8'b10100101;
DRAM[27242] = 8'b10011101;
DRAM[27243] = 8'b10100001;
DRAM[27244] = 8'b10010100;
DRAM[27245] = 8'b1110111;
DRAM[27246] = 8'b1101000;
DRAM[27247] = 8'b1011011;
DRAM[27248] = 8'b1010011;
DRAM[27249] = 8'b1101000;
DRAM[27250] = 8'b10000011;
DRAM[27251] = 8'b1111110;
DRAM[27252] = 8'b1100011;
DRAM[27253] = 8'b1100110;
DRAM[27254] = 8'b1111000;
DRAM[27255] = 8'b1110101;
DRAM[27256] = 8'b1110011;
DRAM[27257] = 8'b10001000;
DRAM[27258] = 8'b10010001;
DRAM[27259] = 8'b10000000;
DRAM[27260] = 8'b10010001;
DRAM[27261] = 8'b10000011;
DRAM[27262] = 8'b10001000;
DRAM[27263] = 8'b10010100;
DRAM[27264] = 8'b10001001;
DRAM[27265] = 8'b10001100;
DRAM[27266] = 8'b10011110;
DRAM[27267] = 8'b10000101;
DRAM[27268] = 8'b10000101;
DRAM[27269] = 8'b10100010;
DRAM[27270] = 8'b10011001;
DRAM[27271] = 8'b10011001;
DRAM[27272] = 8'b10010110;
DRAM[27273] = 8'b10100111;
DRAM[27274] = 8'b10101010;
DRAM[27275] = 8'b10101000;
DRAM[27276] = 8'b10110000;
DRAM[27277] = 8'b10110101;
DRAM[27278] = 8'b10101011;
DRAM[27279] = 8'b10100001;
DRAM[27280] = 8'b10100100;
DRAM[27281] = 8'b10101001;
DRAM[27282] = 8'b10100010;
DRAM[27283] = 8'b10110001;
DRAM[27284] = 8'b10011010;
DRAM[27285] = 8'b10011011;
DRAM[27286] = 8'b10001001;
DRAM[27287] = 8'b10001011;
DRAM[27288] = 8'b10010111;
DRAM[27289] = 8'b10001111;
DRAM[27290] = 8'b10000011;
DRAM[27291] = 8'b10000010;
DRAM[27292] = 8'b10000011;
DRAM[27293] = 8'b1110111;
DRAM[27294] = 8'b1101010;
DRAM[27295] = 8'b1101011;
DRAM[27296] = 8'b1100100;
DRAM[27297] = 8'b1010100;
DRAM[27298] = 8'b1010001;
DRAM[27299] = 8'b1010111;
DRAM[27300] = 8'b1001001;
DRAM[27301] = 8'b100110;
DRAM[27302] = 8'b1111;
DRAM[27303] = 8'b1111;
DRAM[27304] = 8'b10;
DRAM[27305] = 8'b0;
DRAM[27306] = 8'b10011;
DRAM[27307] = 8'b0;
DRAM[27308] = 8'b0;
DRAM[27309] = 8'b11000;
DRAM[27310] = 8'b11001;
DRAM[27311] = 8'b101011;
DRAM[27312] = 8'b1110110;
DRAM[27313] = 8'b10001011;
DRAM[27314] = 8'b10110000;
DRAM[27315] = 8'b11010111;
DRAM[27316] = 8'b11010011;
DRAM[27317] = 8'b11000100;
DRAM[27318] = 8'b11000001;
DRAM[27319] = 8'b10100110;
DRAM[27320] = 8'b10101000;
DRAM[27321] = 8'b10110000;
DRAM[27322] = 8'b10111010;
DRAM[27323] = 8'b11000001;
DRAM[27324] = 8'b11000100;
DRAM[27325] = 8'b10111101;
DRAM[27326] = 8'b10101001;
DRAM[27327] = 8'b10010101;
DRAM[27328] = 8'b10010011;
DRAM[27329] = 8'b10010000;
DRAM[27330] = 8'b10001000;
DRAM[27331] = 8'b1110100;
DRAM[27332] = 8'b1101011;
DRAM[27333] = 8'b1010101;
DRAM[27334] = 8'b1000000;
DRAM[27335] = 8'b1011100;
DRAM[27336] = 8'b10000010;
DRAM[27337] = 8'b10001101;
DRAM[27338] = 8'b10101100;
DRAM[27339] = 8'b10010101;
DRAM[27340] = 8'b10110111;
DRAM[27341] = 8'b11111000;
DRAM[27342] = 8'b11101011;
DRAM[27343] = 8'b11110100;
DRAM[27344] = 8'b11111111;
DRAM[27345] = 8'b11100110;
DRAM[27346] = 8'b11101010;
DRAM[27347] = 8'b11100101;
DRAM[27348] = 8'b11010101;
DRAM[27349] = 8'b11000100;
DRAM[27350] = 8'b10111101;
DRAM[27351] = 8'b11000100;
DRAM[27352] = 8'b10110111;
DRAM[27353] = 8'b10010010;
DRAM[27354] = 8'b10011101;
DRAM[27355] = 8'b10011001;
DRAM[27356] = 8'b10101001;
DRAM[27357] = 8'b10001110;
DRAM[27358] = 8'b10001001;
DRAM[27359] = 8'b10010100;
DRAM[27360] = 8'b10010111;
DRAM[27361] = 8'b10100010;
DRAM[27362] = 8'b10100100;
DRAM[27363] = 8'b11000000;
DRAM[27364] = 8'b11000111;
DRAM[27365] = 8'b10101000;
DRAM[27366] = 8'b10100101;
DRAM[27367] = 8'b10010011;
DRAM[27368] = 8'b10000100;
DRAM[27369] = 8'b1111010;
DRAM[27370] = 8'b1110010;
DRAM[27371] = 8'b1110011;
DRAM[27372] = 8'b1110110;
DRAM[27373] = 8'b1110111;
DRAM[27374] = 8'b1110110;
DRAM[27375] = 8'b1110111;
DRAM[27376] = 8'b1110100;
DRAM[27377] = 8'b1110010;
DRAM[27378] = 8'b1110001;
DRAM[27379] = 8'b1110001;
DRAM[27380] = 8'b1110010;
DRAM[27381] = 8'b1110010;
DRAM[27382] = 8'b1110001;
DRAM[27383] = 8'b1101111;
DRAM[27384] = 8'b1110000;
DRAM[27385] = 8'b1110000;
DRAM[27386] = 8'b1110000;
DRAM[27387] = 8'b1101111;
DRAM[27388] = 8'b1101110;
DRAM[27389] = 8'b1101101;
DRAM[27390] = 8'b1101101;
DRAM[27391] = 8'b1101100;
DRAM[27392] = 8'b10000001;
DRAM[27393] = 8'b10000001;
DRAM[27394] = 8'b10000001;
DRAM[27395] = 8'b10000010;
DRAM[27396] = 8'b10000010;
DRAM[27397] = 8'b10000010;
DRAM[27398] = 8'b10000011;
DRAM[27399] = 8'b10000011;
DRAM[27400] = 8'b10000110;
DRAM[27401] = 8'b10000110;
DRAM[27402] = 8'b10000111;
DRAM[27403] = 8'b10000111;
DRAM[27404] = 8'b10000111;
DRAM[27405] = 8'b10000111;
DRAM[27406] = 8'b10001000;
DRAM[27407] = 8'b10001000;
DRAM[27408] = 8'b10001001;
DRAM[27409] = 8'b10001001;
DRAM[27410] = 8'b10001001;
DRAM[27411] = 8'b10001010;
DRAM[27412] = 8'b10001010;
DRAM[27413] = 8'b10001011;
DRAM[27414] = 8'b10001011;
DRAM[27415] = 8'b10001011;
DRAM[27416] = 8'b10001000;
DRAM[27417] = 8'b10010010;
DRAM[27418] = 8'b10010111;
DRAM[27419] = 8'b10010010;
DRAM[27420] = 8'b10001111;
DRAM[27421] = 8'b10011000;
DRAM[27422] = 8'b10100111;
DRAM[27423] = 8'b10110001;
DRAM[27424] = 8'b10110000;
DRAM[27425] = 8'b11001111;
DRAM[27426] = 8'b11010010;
DRAM[27427] = 8'b10111000;
DRAM[27428] = 8'b10101100;
DRAM[27429] = 8'b10110101;
DRAM[27430] = 8'b10110011;
DRAM[27431] = 8'b10011010;
DRAM[27432] = 8'b10101010;
DRAM[27433] = 8'b10011000;
DRAM[27434] = 8'b10011000;
DRAM[27435] = 8'b10110010;
DRAM[27436] = 8'b10100011;
DRAM[27437] = 8'b10010010;
DRAM[27438] = 8'b10001110;
DRAM[27439] = 8'b10110000;
DRAM[27440] = 8'b10110001;
DRAM[27441] = 8'b10011111;
DRAM[27442] = 8'b10100111;
DRAM[27443] = 8'b10100001;
DRAM[27444] = 8'b10101100;
DRAM[27445] = 8'b10100110;
DRAM[27446] = 8'b10111011;
DRAM[27447] = 8'b10111010;
DRAM[27448] = 8'b11000101;
DRAM[27449] = 8'b10111110;
DRAM[27450] = 8'b11000111;
DRAM[27451] = 8'b11001110;
DRAM[27452] = 8'b11011110;
DRAM[27453] = 8'b11001110;
DRAM[27454] = 8'b11100001;
DRAM[27455] = 8'b11011001;
DRAM[27456] = 8'b11010100;
DRAM[27457] = 8'b11010101;
DRAM[27458] = 8'b11011011;
DRAM[27459] = 8'b11011011;
DRAM[27460] = 8'b11100011;
DRAM[27461] = 8'b11010100;
DRAM[27462] = 8'b10110000;
DRAM[27463] = 8'b10010100;
DRAM[27464] = 8'b10110001;
DRAM[27465] = 8'b10000110;
DRAM[27466] = 8'b1000111;
DRAM[27467] = 8'b1001000;
DRAM[27468] = 8'b1010010;
DRAM[27469] = 8'b1100101;
DRAM[27470] = 8'b1100100;
DRAM[27471] = 8'b1111111;
DRAM[27472] = 8'b10010110;
DRAM[27473] = 8'b10100000;
DRAM[27474] = 8'b10100111;
DRAM[27475] = 8'b10110101;
DRAM[27476] = 8'b11001011;
DRAM[27477] = 8'b11001110;
DRAM[27478] = 8'b11000100;
DRAM[27479] = 8'b11000010;
DRAM[27480] = 8'b11000110;
DRAM[27481] = 8'b11010001;
DRAM[27482] = 8'b11011011;
DRAM[27483] = 8'b11011011;
DRAM[27484] = 8'b11011001;
DRAM[27485] = 8'b11011011;
DRAM[27486] = 8'b11100010;
DRAM[27487] = 8'b11101001;
DRAM[27488] = 8'b11101000;
DRAM[27489] = 8'b11011100;
DRAM[27490] = 8'b11001111;
DRAM[27491] = 8'b11001101;
DRAM[27492] = 8'b11010011;
DRAM[27493] = 8'b11010001;
DRAM[27494] = 8'b11000000;
DRAM[27495] = 8'b10101110;
DRAM[27496] = 8'b10011111;
DRAM[27497] = 8'b10011001;
DRAM[27498] = 8'b1111111;
DRAM[27499] = 8'b10001101;
DRAM[27500] = 8'b10001100;
DRAM[27501] = 8'b1110100;
DRAM[27502] = 8'b1110101;
DRAM[27503] = 8'b1100110;
DRAM[27504] = 8'b1100010;
DRAM[27505] = 8'b1011010;
DRAM[27506] = 8'b1101110;
DRAM[27507] = 8'b1110111;
DRAM[27508] = 8'b1100110;
DRAM[27509] = 8'b1101111;
DRAM[27510] = 8'b1111111;
DRAM[27511] = 8'b1110011;
DRAM[27512] = 8'b1110101;
DRAM[27513] = 8'b10000010;
DRAM[27514] = 8'b10001100;
DRAM[27515] = 8'b1111111;
DRAM[27516] = 8'b10001110;
DRAM[27517] = 8'b1111111;
DRAM[27518] = 8'b10000011;
DRAM[27519] = 8'b10001010;
DRAM[27520] = 8'b10001011;
DRAM[27521] = 8'b10010010;
DRAM[27522] = 8'b10010101;
DRAM[27523] = 8'b1111101;
DRAM[27524] = 8'b10000110;
DRAM[27525] = 8'b10100000;
DRAM[27526] = 8'b10011010;
DRAM[27527] = 8'b10100000;
DRAM[27528] = 8'b10011100;
DRAM[27529] = 8'b10110000;
DRAM[27530] = 8'b10101100;
DRAM[27531] = 8'b10100010;
DRAM[27532] = 8'b10101100;
DRAM[27533] = 8'b10101111;
DRAM[27534] = 8'b10101010;
DRAM[27535] = 8'b10110000;
DRAM[27536] = 8'b10011111;
DRAM[27537] = 8'b10101111;
DRAM[27538] = 8'b10101010;
DRAM[27539] = 8'b10101101;
DRAM[27540] = 8'b10100100;
DRAM[27541] = 8'b10100010;
DRAM[27542] = 8'b10001110;
DRAM[27543] = 8'b10001110;
DRAM[27544] = 8'b10001001;
DRAM[27545] = 8'b10001110;
DRAM[27546] = 8'b10000001;
DRAM[27547] = 8'b1111011;
DRAM[27548] = 8'b10000011;
DRAM[27549] = 8'b1110111;
DRAM[27550] = 8'b1101000;
DRAM[27551] = 8'b1101111;
DRAM[27552] = 8'b1011101;
DRAM[27553] = 8'b1001101;
DRAM[27554] = 8'b1001010;
DRAM[27555] = 8'b1010011;
DRAM[27556] = 8'b1000011;
DRAM[27557] = 8'b11100;
DRAM[27558] = 8'b101;
DRAM[27559] = 8'b111;
DRAM[27560] = 8'b1001;
DRAM[27561] = 8'b11111;
DRAM[27562] = 8'b11010;
DRAM[27563] = 8'b1110;
DRAM[27564] = 8'b10101;
DRAM[27565] = 8'b10000;
DRAM[27566] = 8'b100;
DRAM[27567] = 8'b100100;
DRAM[27568] = 8'b0;
DRAM[27569] = 8'b11001;
DRAM[27570] = 8'b1010001;
DRAM[27571] = 8'b1111101;
DRAM[27572] = 8'b10101010;
DRAM[27573] = 8'b11100011;
DRAM[27574] = 8'b11010111;
DRAM[27575] = 8'b10000000;
DRAM[27576] = 8'b1111100;
DRAM[27577] = 8'b10011000;
DRAM[27578] = 8'b10101111;
DRAM[27579] = 8'b10110011;
DRAM[27580] = 8'b10110001;
DRAM[27581] = 8'b10110011;
DRAM[27582] = 8'b10110000;
DRAM[27583] = 8'b10101000;
DRAM[27584] = 8'b10001111;
DRAM[27585] = 8'b10000111;
DRAM[27586] = 8'b10000001;
DRAM[27587] = 8'b1110000;
DRAM[27588] = 8'b1100110;
DRAM[27589] = 8'b1010010;
DRAM[27590] = 8'b111010;
DRAM[27591] = 8'b1001010;
DRAM[27592] = 8'b1110111;
DRAM[27593] = 8'b1111110;
DRAM[27594] = 8'b10011011;
DRAM[27595] = 8'b10011000;
DRAM[27596] = 8'b10110111;
DRAM[27597] = 8'b11100100;
DRAM[27598] = 8'b11100010;
DRAM[27599] = 8'b11111000;
DRAM[27600] = 8'b11111011;
DRAM[27601] = 8'b11100110;
DRAM[27602] = 8'b11101100;
DRAM[27603] = 8'b11101101;
DRAM[27604] = 8'b11010011;
DRAM[27605] = 8'b11010011;
DRAM[27606] = 8'b10101110;
DRAM[27607] = 8'b10110000;
DRAM[27608] = 8'b10111011;
DRAM[27609] = 8'b10010101;
DRAM[27610] = 8'b10011001;
DRAM[27611] = 8'b10011010;
DRAM[27612] = 8'b10100101;
DRAM[27613] = 8'b10010010;
DRAM[27614] = 8'b10001001;
DRAM[27615] = 8'b10010110;
DRAM[27616] = 8'b10011111;
DRAM[27617] = 8'b10101111;
DRAM[27618] = 8'b10101110;
DRAM[27619] = 8'b11000111;
DRAM[27620] = 8'b11000110;
DRAM[27621] = 8'b10010100;
DRAM[27622] = 8'b10011101;
DRAM[27623] = 8'b10000011;
DRAM[27624] = 8'b10000100;
DRAM[27625] = 8'b1111011;
DRAM[27626] = 8'b1110110;
DRAM[27627] = 8'b1110111;
DRAM[27628] = 8'b1111001;
DRAM[27629] = 8'b1110110;
DRAM[27630] = 8'b1110100;
DRAM[27631] = 8'b1110100;
DRAM[27632] = 8'b1110100;
DRAM[27633] = 8'b1110010;
DRAM[27634] = 8'b1110001;
DRAM[27635] = 8'b1110001;
DRAM[27636] = 8'b1110010;
DRAM[27637] = 8'b1110011;
DRAM[27638] = 8'b1110001;
DRAM[27639] = 8'b1110000;
DRAM[27640] = 8'b1110001;
DRAM[27641] = 8'b1110001;
DRAM[27642] = 8'b1110000;
DRAM[27643] = 8'b1101111;
DRAM[27644] = 8'b1101110;
DRAM[27645] = 8'b1101110;
DRAM[27646] = 8'b1101101;
DRAM[27647] = 8'b1101101;
DRAM[27648] = 8'b10000011;
DRAM[27649] = 8'b10000011;
DRAM[27650] = 8'b10000011;
DRAM[27651] = 8'b10000100;
DRAM[27652] = 8'b10000100;
DRAM[27653] = 8'b10000101;
DRAM[27654] = 8'b10000101;
DRAM[27655] = 8'b10000101;
DRAM[27656] = 8'b10000110;
DRAM[27657] = 8'b10000110;
DRAM[27658] = 8'b10000111;
DRAM[27659] = 8'b10000111;
DRAM[27660] = 8'b10001000;
DRAM[27661] = 8'b10001000;
DRAM[27662] = 8'b10001000;
DRAM[27663] = 8'b10001001;
DRAM[27664] = 8'b10001001;
DRAM[27665] = 8'b10001001;
DRAM[27666] = 8'b10001010;
DRAM[27667] = 8'b10001010;
DRAM[27668] = 8'b10001011;
DRAM[27669] = 8'b10001011;
DRAM[27670] = 8'b10001011;
DRAM[27671] = 8'b10001011;
DRAM[27672] = 8'b10001011;
DRAM[27673] = 8'b10001111;
DRAM[27674] = 8'b10001110;
DRAM[27675] = 8'b10001000;
DRAM[27676] = 8'b10001001;
DRAM[27677] = 8'b10010101;
DRAM[27678] = 8'b10100011;
DRAM[27679] = 8'b10101010;
DRAM[27680] = 8'b10110011;
DRAM[27681] = 8'b11000001;
DRAM[27682] = 8'b11010000;
DRAM[27683] = 8'b11001001;
DRAM[27684] = 8'b10111011;
DRAM[27685] = 8'b10110001;
DRAM[27686] = 8'b10101001;
DRAM[27687] = 8'b10101001;
DRAM[27688] = 8'b10100000;
DRAM[27689] = 8'b10011001;
DRAM[27690] = 8'b10100010;
DRAM[27691] = 8'b10100011;
DRAM[27692] = 8'b10011101;
DRAM[27693] = 8'b10000010;
DRAM[27694] = 8'b10010110;
DRAM[27695] = 8'b10101110;
DRAM[27696] = 8'b10100110;
DRAM[27697] = 8'b10011010;
DRAM[27698] = 8'b10101000;
DRAM[27699] = 8'b10100010;
DRAM[27700] = 8'b10101100;
DRAM[27701] = 8'b10100111;
DRAM[27702] = 8'b10111010;
DRAM[27703] = 8'b10111000;
DRAM[27704] = 8'b11001011;
DRAM[27705] = 8'b10111110;
DRAM[27706] = 8'b11001011;
DRAM[27707] = 8'b11010110;
DRAM[27708] = 8'b11100001;
DRAM[27709] = 8'b11010001;
DRAM[27710] = 8'b11101000;
DRAM[27711] = 8'b11011101;
DRAM[27712] = 8'b11010000;
DRAM[27713] = 8'b11010111;
DRAM[27714] = 8'b11011011;
DRAM[27715] = 8'b11100110;
DRAM[27716] = 8'b11011101;
DRAM[27717] = 8'b11001100;
DRAM[27718] = 8'b10101110;
DRAM[27719] = 8'b10010010;
DRAM[27720] = 8'b10110101;
DRAM[27721] = 8'b10000000;
DRAM[27722] = 8'b1000101;
DRAM[27723] = 8'b1010001;
DRAM[27724] = 8'b1011001;
DRAM[27725] = 8'b1101010;
DRAM[27726] = 8'b1101011;
DRAM[27727] = 8'b10000101;
DRAM[27728] = 8'b10001101;
DRAM[27729] = 8'b10011101;
DRAM[27730] = 8'b10100100;
DRAM[27731] = 8'b10100111;
DRAM[27732] = 8'b10101110;
DRAM[27733] = 8'b10110101;
DRAM[27734] = 8'b11000010;
DRAM[27735] = 8'b11010110;
DRAM[27736] = 8'b11001001;
DRAM[27737] = 8'b11011110;
DRAM[27738] = 8'b11101000;
DRAM[27739] = 8'b11011111;
DRAM[27740] = 8'b11011110;
DRAM[27741] = 8'b11101011;
DRAM[27742] = 8'b11110001;
DRAM[27743] = 8'b11101101;
DRAM[27744] = 8'b11010100;
DRAM[27745] = 8'b11000100;
DRAM[27746] = 8'b10111000;
DRAM[27747] = 8'b10110101;
DRAM[27748] = 8'b10101110;
DRAM[27749] = 8'b10100110;
DRAM[27750] = 8'b10101011;
DRAM[27751] = 8'b10111001;
DRAM[27752] = 8'b10011100;
DRAM[27753] = 8'b10010000;
DRAM[27754] = 8'b1110000;
DRAM[27755] = 8'b1111100;
DRAM[27756] = 8'b10000011;
DRAM[27757] = 8'b1110011;
DRAM[27758] = 8'b1110110;
DRAM[27759] = 8'b1100011;
DRAM[27760] = 8'b1110000;
DRAM[27761] = 8'b1010010;
DRAM[27762] = 8'b1011110;
DRAM[27763] = 8'b1110100;
DRAM[27764] = 8'b1100111;
DRAM[27765] = 8'b1100001;
DRAM[27766] = 8'b1101010;
DRAM[27767] = 8'b1100100;
DRAM[27768] = 8'b1110101;
DRAM[27769] = 8'b1111000;
DRAM[27770] = 8'b10000101;
DRAM[27771] = 8'b10000000;
DRAM[27772] = 8'b10010001;
DRAM[27773] = 8'b10000100;
DRAM[27774] = 8'b10000110;
DRAM[27775] = 8'b10000011;
DRAM[27776] = 8'b10010010;
DRAM[27777] = 8'b10010010;
DRAM[27778] = 8'b10010011;
DRAM[27779] = 8'b10001101;
DRAM[27780] = 8'b10010110;
DRAM[27781] = 8'b10011111;
DRAM[27782] = 8'b10011101;
DRAM[27783] = 8'b10101010;
DRAM[27784] = 8'b10100001;
DRAM[27785] = 8'b10110100;
DRAM[27786] = 8'b10101111;
DRAM[27787] = 8'b10100101;
DRAM[27788] = 8'b10101101;
DRAM[27789] = 8'b10101110;
DRAM[27790] = 8'b10101001;
DRAM[27791] = 8'b10110010;
DRAM[27792] = 8'b10101111;
DRAM[27793] = 8'b10110111;
DRAM[27794] = 8'b10111010;
DRAM[27795] = 8'b10100111;
DRAM[27796] = 8'b10101011;
DRAM[27797] = 8'b10011010;
DRAM[27798] = 8'b10010011;
DRAM[27799] = 8'b10001011;
DRAM[27800] = 8'b10001001;
DRAM[27801] = 8'b10010100;
DRAM[27802] = 8'b10001010;
DRAM[27803] = 8'b10000001;
DRAM[27804] = 8'b10001000;
DRAM[27805] = 8'b1111111;
DRAM[27806] = 8'b1110000;
DRAM[27807] = 8'b1110100;
DRAM[27808] = 8'b1100010;
DRAM[27809] = 8'b1001100;
DRAM[27810] = 8'b1000001;
DRAM[27811] = 8'b1000010;
DRAM[27812] = 8'b110010;
DRAM[27813] = 8'b10001;
DRAM[27814] = 8'b0;
DRAM[27815] = 8'b100;
DRAM[27816] = 8'b11111;
DRAM[27817] = 8'b11111;
DRAM[27818] = 8'b1100;
DRAM[27819] = 8'b111001;
DRAM[27820] = 8'b111;
DRAM[27821] = 8'b0;
DRAM[27822] = 8'b10011;
DRAM[27823] = 8'b10000;
DRAM[27824] = 8'b101010;
DRAM[27825] = 8'b10001;
DRAM[27826] = 8'b10100;
DRAM[27827] = 8'b11010;
DRAM[27828] = 8'b101010;
DRAM[27829] = 8'b1110000;
DRAM[27830] = 8'b10110111;
DRAM[27831] = 8'b11001100;
DRAM[27832] = 8'b10001010;
DRAM[27833] = 8'b10000111;
DRAM[27834] = 8'b10010111;
DRAM[27835] = 8'b10110000;
DRAM[27836] = 8'b10110001;
DRAM[27837] = 8'b10011110;
DRAM[27838] = 8'b10011101;
DRAM[27839] = 8'b10101101;
DRAM[27840] = 8'b10010100;
DRAM[27841] = 8'b10000110;
DRAM[27842] = 8'b10000001;
DRAM[27843] = 8'b1110000;
DRAM[27844] = 8'b1100011;
DRAM[27845] = 8'b1010100;
DRAM[27846] = 8'b111111;
DRAM[27847] = 8'b1001000;
DRAM[27848] = 8'b1011111;
DRAM[27849] = 8'b1111010;
DRAM[27850] = 8'b10001100;
DRAM[27851] = 8'b10011101;
DRAM[27852] = 8'b10111010;
DRAM[27853] = 8'b11010011;
DRAM[27854] = 8'b11100100;
DRAM[27855] = 8'b11101111;
DRAM[27856] = 8'b11111011;
DRAM[27857] = 8'b11110000;
DRAM[27858] = 8'b11110001;
DRAM[27859] = 8'b11101110;
DRAM[27860] = 8'b11010010;
DRAM[27861] = 8'b11100001;
DRAM[27862] = 8'b10101111;
DRAM[27863] = 8'b10011110;
DRAM[27864] = 8'b10110111;
DRAM[27865] = 8'b10100001;
DRAM[27866] = 8'b10010110;
DRAM[27867] = 8'b10011011;
DRAM[27868] = 8'b10010101;
DRAM[27869] = 8'b10011101;
DRAM[27870] = 8'b10001010;
DRAM[27871] = 8'b10010101;
DRAM[27872] = 8'b10100011;
DRAM[27873] = 8'b10111000;
DRAM[27874] = 8'b10110101;
DRAM[27875] = 8'b10111111;
DRAM[27876] = 8'b11000001;
DRAM[27877] = 8'b10001001;
DRAM[27878] = 8'b10010101;
DRAM[27879] = 8'b1111100;
DRAM[27880] = 8'b10000000;
DRAM[27881] = 8'b1111001;
DRAM[27882] = 8'b1110110;
DRAM[27883] = 8'b1111000;
DRAM[27884] = 8'b1111001;
DRAM[27885] = 8'b1110110;
DRAM[27886] = 8'b1110100;
DRAM[27887] = 8'b1110100;
DRAM[27888] = 8'b1110100;
DRAM[27889] = 8'b1110011;
DRAM[27890] = 8'b1110001;
DRAM[27891] = 8'b1110010;
DRAM[27892] = 8'b1110011;
DRAM[27893] = 8'b1110011;
DRAM[27894] = 8'b1110010;
DRAM[27895] = 8'b1110000;
DRAM[27896] = 8'b1110001;
DRAM[27897] = 8'b1110001;
DRAM[27898] = 8'b1110000;
DRAM[27899] = 8'b1110000;
DRAM[27900] = 8'b1101111;
DRAM[27901] = 8'b1101110;
DRAM[27902] = 8'b1101101;
DRAM[27903] = 8'b1101101;
DRAM[27904] = 8'b10000101;
DRAM[27905] = 8'b10000101;
DRAM[27906] = 8'b10000101;
DRAM[27907] = 8'b10000110;
DRAM[27908] = 8'b10000110;
DRAM[27909] = 8'b10000110;
DRAM[27910] = 8'b10000111;
DRAM[27911] = 8'b10000111;
DRAM[27912] = 8'b10000101;
DRAM[27913] = 8'b10000101;
DRAM[27914] = 8'b10000110;
DRAM[27915] = 8'b10000111;
DRAM[27916] = 8'b10000111;
DRAM[27917] = 8'b10001000;
DRAM[27918] = 8'b10001001;
DRAM[27919] = 8'b10001001;
DRAM[27920] = 8'b10001001;
DRAM[27921] = 8'b10001001;
DRAM[27922] = 8'b10001001;
DRAM[27923] = 8'b10001010;
DRAM[27924] = 8'b10001010;
DRAM[27925] = 8'b10001011;
DRAM[27926] = 8'b10001011;
DRAM[27927] = 8'b10001011;
DRAM[27928] = 8'b10001110;
DRAM[27929] = 8'b10001010;
DRAM[27930] = 8'b10000110;
DRAM[27931] = 8'b10000110;
DRAM[27932] = 8'b10001010;
DRAM[27933] = 8'b10010011;
DRAM[27934] = 8'b10011110;
DRAM[27935] = 8'b10100110;
DRAM[27936] = 8'b10110100;
DRAM[27937] = 8'b10110100;
DRAM[27938] = 8'b11001010;
DRAM[27939] = 8'b11001111;
DRAM[27940] = 8'b11000011;
DRAM[27941] = 8'b10110010;
DRAM[27942] = 8'b10100011;
DRAM[27943] = 8'b10110001;
DRAM[27944] = 8'b10011001;
DRAM[27945] = 8'b10011100;
DRAM[27946] = 8'b10100001;
DRAM[27947] = 8'b10010100;
DRAM[27948] = 8'b10010101;
DRAM[27949] = 8'b1111100;
DRAM[27950] = 8'b10011100;
DRAM[27951] = 8'b10100110;
DRAM[27952] = 8'b10011110;
DRAM[27953] = 8'b10100001;
DRAM[27954] = 8'b10100111;
DRAM[27955] = 8'b10100001;
DRAM[27956] = 8'b10100110;
DRAM[27957] = 8'b10100011;
DRAM[27958] = 8'b10101110;
DRAM[27959] = 8'b10110110;
DRAM[27960] = 8'b11001101;
DRAM[27961] = 8'b10111011;
DRAM[27962] = 8'b11010000;
DRAM[27963] = 8'b11011011;
DRAM[27964] = 8'b11011011;
DRAM[27965] = 8'b11011100;
DRAM[27966] = 8'b11100110;
DRAM[27967] = 8'b11011110;
DRAM[27968] = 8'b11101001;
DRAM[27969] = 8'b11011001;
DRAM[27970] = 8'b11010000;
DRAM[27971] = 8'b11101101;
DRAM[27972] = 8'b11010111;
DRAM[27973] = 8'b10111001;
DRAM[27974] = 8'b10101010;
DRAM[27975] = 8'b10100011;
DRAM[27976] = 8'b10100011;
DRAM[27977] = 8'b1101111;
DRAM[27978] = 8'b1001001;
DRAM[27979] = 8'b1011001;
DRAM[27980] = 8'b1100111;
DRAM[27981] = 8'b1101111;
DRAM[27982] = 8'b1110011;
DRAM[27983] = 8'b10000100;
DRAM[27984] = 8'b10001010;
DRAM[27985] = 8'b10011001;
DRAM[27986] = 8'b10100010;
DRAM[27987] = 8'b10101011;
DRAM[27988] = 8'b10111010;
DRAM[27989] = 8'b11000011;
DRAM[27990] = 8'b11001101;
DRAM[27991] = 8'b11011101;
DRAM[27992] = 8'b11010010;
DRAM[27993] = 8'b11011010;
DRAM[27994] = 8'b11011001;
DRAM[27995] = 8'b11010100;
DRAM[27996] = 8'b11011110;
DRAM[27997] = 8'b11101100;
DRAM[27998] = 8'b11100110;
DRAM[27999] = 8'b11010010;
DRAM[28000] = 8'b11000011;
DRAM[28001] = 8'b10110110;
DRAM[28002] = 8'b10110000;
DRAM[28003] = 8'b10110101;
DRAM[28004] = 8'b10110001;
DRAM[28005] = 8'b10100011;
DRAM[28006] = 8'b10011011;
DRAM[28007] = 8'b10011110;
DRAM[28008] = 8'b10001011;
DRAM[28009] = 8'b10000010;
DRAM[28010] = 8'b1101110;
DRAM[28011] = 8'b1110000;
DRAM[28012] = 8'b1110010;
DRAM[28013] = 8'b1100110;
DRAM[28014] = 8'b1011001;
DRAM[28015] = 8'b1000010;
DRAM[28016] = 8'b1011000;
DRAM[28017] = 8'b1000100;
DRAM[28018] = 8'b1010111;
DRAM[28019] = 8'b1110101;
DRAM[28020] = 8'b1101000;
DRAM[28021] = 8'b1010100;
DRAM[28022] = 8'b1011001;
DRAM[28023] = 8'b1100100;
DRAM[28024] = 8'b1101111;
DRAM[28025] = 8'b1101100;
DRAM[28026] = 8'b1111100;
DRAM[28027] = 8'b10000000;
DRAM[28028] = 8'b10010010;
DRAM[28029] = 8'b10001000;
DRAM[28030] = 8'b10001101;
DRAM[28031] = 8'b10000110;
DRAM[28032] = 8'b10001110;
DRAM[28033] = 8'b10001001;
DRAM[28034] = 8'b10010001;
DRAM[28035] = 8'b10011111;
DRAM[28036] = 8'b10100000;
DRAM[28037] = 8'b10011011;
DRAM[28038] = 8'b10011110;
DRAM[28039] = 8'b10101000;
DRAM[28040] = 8'b10100100;
DRAM[28041] = 8'b10110000;
DRAM[28042] = 8'b10110011;
DRAM[28043] = 8'b10110010;
DRAM[28044] = 8'b10110110;
DRAM[28045] = 8'b10110100;
DRAM[28046] = 8'b10101100;
DRAM[28047] = 8'b10101010;
DRAM[28048] = 8'b10110110;
DRAM[28049] = 8'b10110010;
DRAM[28050] = 8'b10111100;
DRAM[28051] = 8'b10100111;
DRAM[28052] = 8'b10101101;
DRAM[28053] = 8'b10011010;
DRAM[28054] = 8'b10100000;
DRAM[28055] = 8'b10010101;
DRAM[28056] = 8'b10010010;
DRAM[28057] = 8'b10011010;
DRAM[28058] = 8'b10010110;
DRAM[28059] = 8'b10001100;
DRAM[28060] = 8'b10001011;
DRAM[28061] = 8'b10000101;
DRAM[28062] = 8'b1110110;
DRAM[28063] = 8'b1101101;
DRAM[28064] = 8'b1101010;
DRAM[28065] = 8'b1001110;
DRAM[28066] = 8'b110100;
DRAM[28067] = 8'b100111;
DRAM[28068] = 8'b11001;
DRAM[28069] = 8'b1000;
DRAM[28070] = 8'b0;
DRAM[28071] = 8'b101;
DRAM[28072] = 8'b10011;
DRAM[28073] = 8'b1111011;
DRAM[28074] = 8'b11001;
DRAM[28075] = 8'b1010;
DRAM[28076] = 8'b10001;
DRAM[28077] = 8'b1101;
DRAM[28078] = 8'b0;
DRAM[28079] = 8'b101;
DRAM[28080] = 8'b10111;
DRAM[28081] = 8'b1011;
DRAM[28082] = 8'b100011;
DRAM[28083] = 8'b100000;
DRAM[28084] = 8'b0;
DRAM[28085] = 8'b100;
DRAM[28086] = 8'b110011;
DRAM[28087] = 8'b1101011;
DRAM[28088] = 8'b10010110;
DRAM[28089] = 8'b10010000;
DRAM[28090] = 8'b10010001;
DRAM[28091] = 8'b10011110;
DRAM[28092] = 8'b10101010;
DRAM[28093] = 8'b10101001;
DRAM[28094] = 8'b10011100;
DRAM[28095] = 8'b10010001;
DRAM[28096] = 8'b10010101;
DRAM[28097] = 8'b10000100;
DRAM[28098] = 8'b1111111;
DRAM[28099] = 8'b1101101;
DRAM[28100] = 8'b1011100;
DRAM[28101] = 8'b1010011;
DRAM[28102] = 8'b1000011;
DRAM[28103] = 8'b1001000;
DRAM[28104] = 8'b1000101;
DRAM[28105] = 8'b1111001;
DRAM[28106] = 8'b10001010;
DRAM[28107] = 8'b10010111;
DRAM[28108] = 8'b10110001;
DRAM[28109] = 8'b11001100;
DRAM[28110] = 8'b11100101;
DRAM[28111] = 8'b11100000;
DRAM[28112] = 8'b11111111;
DRAM[28113] = 8'b11111100;
DRAM[28114] = 8'b11110100;
DRAM[28115] = 8'b11101110;
DRAM[28116] = 8'b11010110;
DRAM[28117] = 8'b11100101;
DRAM[28118] = 8'b11000001;
DRAM[28119] = 8'b10100100;
DRAM[28120] = 8'b10110010;
DRAM[28121] = 8'b10100110;
DRAM[28122] = 8'b10010110;
DRAM[28123] = 8'b10010111;
DRAM[28124] = 8'b10001010;
DRAM[28125] = 8'b10100001;
DRAM[28126] = 8'b10001101;
DRAM[28127] = 8'b10010110;
DRAM[28128] = 8'b10100000;
DRAM[28129] = 8'b10111100;
DRAM[28130] = 8'b10111000;
DRAM[28131] = 8'b10100111;
DRAM[28132] = 8'b10111000;
DRAM[28133] = 8'b10000111;
DRAM[28134] = 8'b10001011;
DRAM[28135] = 8'b1111110;
DRAM[28136] = 8'b1111001;
DRAM[28137] = 8'b1110100;
DRAM[28138] = 8'b1110010;
DRAM[28139] = 8'b1110101;
DRAM[28140] = 8'b1110111;
DRAM[28141] = 8'b1110101;
DRAM[28142] = 8'b1110100;
DRAM[28143] = 8'b1110110;
DRAM[28144] = 8'b1110101;
DRAM[28145] = 8'b1110011;
DRAM[28146] = 8'b1110010;
DRAM[28147] = 8'b1110010;
DRAM[28148] = 8'b1110011;
DRAM[28149] = 8'b1110011;
DRAM[28150] = 8'b1110010;
DRAM[28151] = 8'b1110000;
DRAM[28152] = 8'b1110010;
DRAM[28153] = 8'b1110001;
DRAM[28154] = 8'b1110001;
DRAM[28155] = 8'b1110000;
DRAM[28156] = 8'b1101111;
DRAM[28157] = 8'b1101110;
DRAM[28158] = 8'b1101110;
DRAM[28159] = 8'b1101110;
DRAM[28160] = 8'b10000101;
DRAM[28161] = 8'b10000110;
DRAM[28162] = 8'b10000110;
DRAM[28163] = 8'b10000110;
DRAM[28164] = 8'b10000111;
DRAM[28165] = 8'b10000111;
DRAM[28166] = 8'b10000111;
DRAM[28167] = 8'b10001000;
DRAM[28168] = 8'b10000100;
DRAM[28169] = 8'b10000100;
DRAM[28170] = 8'b10000101;
DRAM[28171] = 8'b10000110;
DRAM[28172] = 8'b10000111;
DRAM[28173] = 8'b10001000;
DRAM[28174] = 8'b10001000;
DRAM[28175] = 8'b10001001;
DRAM[28176] = 8'b10001000;
DRAM[28177] = 8'b10001001;
DRAM[28178] = 8'b10001001;
DRAM[28179] = 8'b10001001;
DRAM[28180] = 8'b10001010;
DRAM[28181] = 8'b10001010;
DRAM[28182] = 8'b10001010;
DRAM[28183] = 8'b10001010;
DRAM[28184] = 8'b10001111;
DRAM[28185] = 8'b10001000;
DRAM[28186] = 8'b10000111;
DRAM[28187] = 8'b10001101;
DRAM[28188] = 8'b10010000;
DRAM[28189] = 8'b10010000;
DRAM[28190] = 8'b10011000;
DRAM[28191] = 8'b10100100;
DRAM[28192] = 8'b10100111;
DRAM[28193] = 8'b10101001;
DRAM[28194] = 8'b11000001;
DRAM[28195] = 8'b11000001;
DRAM[28196] = 8'b11000000;
DRAM[28197] = 8'b11000001;
DRAM[28198] = 8'b10101101;
DRAM[28199] = 8'b10110000;
DRAM[28200] = 8'b10011110;
DRAM[28201] = 8'b10100010;
DRAM[28202] = 8'b10010101;
DRAM[28203] = 8'b10010100;
DRAM[28204] = 8'b10010000;
DRAM[28205] = 8'b10000101;
DRAM[28206] = 8'b10011110;
DRAM[28207] = 8'b10100010;
DRAM[28208] = 8'b10011011;
DRAM[28209] = 8'b10101101;
DRAM[28210] = 8'b10100100;
DRAM[28211] = 8'b10011111;
DRAM[28212] = 8'b10011110;
DRAM[28213] = 8'b10100001;
DRAM[28214] = 8'b10100011;
DRAM[28215] = 8'b10111011;
DRAM[28216] = 8'b11001100;
DRAM[28217] = 8'b10110111;
DRAM[28218] = 8'b11010011;
DRAM[28219] = 8'b11011101;
DRAM[28220] = 8'b11001111;
DRAM[28221] = 8'b11100110;
DRAM[28222] = 8'b11011101;
DRAM[28223] = 8'b11011010;
DRAM[28224] = 8'b11110100;
DRAM[28225] = 8'b11011100;
DRAM[28226] = 8'b11000100;
DRAM[28227] = 8'b11100101;
DRAM[28228] = 8'b11001010;
DRAM[28229] = 8'b10110011;
DRAM[28230] = 8'b10101110;
DRAM[28231] = 8'b10101000;
DRAM[28232] = 8'b10010011;
DRAM[28233] = 8'b1100001;
DRAM[28234] = 8'b1001100;
DRAM[28235] = 8'b1010110;
DRAM[28236] = 8'b1101001;
DRAM[28237] = 8'b1101000;
DRAM[28238] = 8'b1110110;
DRAM[28239] = 8'b10000000;
DRAM[28240] = 8'b10010000;
DRAM[28241] = 8'b10011101;
DRAM[28242] = 8'b10101000;
DRAM[28243] = 8'b10111000;
DRAM[28244] = 8'b11001110;
DRAM[28245] = 8'b11010011;
DRAM[28246] = 8'b11001111;
DRAM[28247] = 8'b11010010;
DRAM[28248] = 8'b11100000;
DRAM[28249] = 8'b11011000;
DRAM[28250] = 8'b11010100;
DRAM[28251] = 8'b11011011;
DRAM[28252] = 8'b11100100;
DRAM[28253] = 8'b11100011;
DRAM[28254] = 8'b11010110;
DRAM[28255] = 8'b11001001;
DRAM[28256] = 8'b11001010;
DRAM[28257] = 8'b11001000;
DRAM[28258] = 8'b11000100;
DRAM[28259] = 8'b11000010;
DRAM[28260] = 8'b11000001;
DRAM[28261] = 8'b10110110;
DRAM[28262] = 8'b10011011;
DRAM[28263] = 8'b10000001;
DRAM[28264] = 8'b1110011;
DRAM[28265] = 8'b1101100;
DRAM[28266] = 8'b1100111;
DRAM[28267] = 8'b1010110;
DRAM[28268] = 8'b1010110;
DRAM[28269] = 8'b1100000;
DRAM[28270] = 8'b1010110;
DRAM[28271] = 8'b1001111;
DRAM[28272] = 8'b111010;
DRAM[28273] = 8'b111000;
DRAM[28274] = 8'b1001100;
DRAM[28275] = 8'b1100111;
DRAM[28276] = 8'b1100111;
DRAM[28277] = 8'b1010111;
DRAM[28278] = 8'b1011010;
DRAM[28279] = 8'b1101011;
DRAM[28280] = 8'b1101001;
DRAM[28281] = 8'b1100011;
DRAM[28282] = 8'b1111000;
DRAM[28283] = 8'b1111110;
DRAM[28284] = 8'b10001100;
DRAM[28285] = 8'b10000100;
DRAM[28286] = 8'b10010000;
DRAM[28287] = 8'b10001011;
DRAM[28288] = 8'b10001110;
DRAM[28289] = 8'b10000100;
DRAM[28290] = 8'b10001111;
DRAM[28291] = 8'b10100001;
DRAM[28292] = 8'b10011000;
DRAM[28293] = 8'b10010100;
DRAM[28294] = 8'b10100101;
DRAM[28295] = 8'b10100111;
DRAM[28296] = 8'b10101100;
DRAM[28297] = 8'b10101100;
DRAM[28298] = 8'b10110011;
DRAM[28299] = 8'b10111010;
DRAM[28300] = 8'b10111001;
DRAM[28301] = 8'b10111011;
DRAM[28302] = 8'b10110111;
DRAM[28303] = 8'b10101001;
DRAM[28304] = 8'b10110110;
DRAM[28305] = 8'b10101010;
DRAM[28306] = 8'b10110010;
DRAM[28307] = 8'b10110010;
DRAM[28308] = 8'b10100111;
DRAM[28309] = 8'b10100011;
DRAM[28310] = 8'b10101100;
DRAM[28311] = 8'b10100100;
DRAM[28312] = 8'b10011010;
DRAM[28313] = 8'b10011100;
DRAM[28314] = 8'b10011110;
DRAM[28315] = 8'b10010110;
DRAM[28316] = 8'b10001100;
DRAM[28317] = 8'b10001010;
DRAM[28318] = 8'b1111101;
DRAM[28319] = 8'b1100101;
DRAM[28320] = 8'b1100100;
DRAM[28321] = 8'b1001010;
DRAM[28322] = 8'b101010;
DRAM[28323] = 8'b10111;
DRAM[28324] = 8'b10000;
DRAM[28325] = 8'b1011;
DRAM[28326] = 8'b1000;
DRAM[28327] = 8'b110;
DRAM[28328] = 8'b10100;
DRAM[28329] = 8'b110110;
DRAM[28330] = 8'b0;
DRAM[28331] = 8'b1011;
DRAM[28332] = 8'b1000;
DRAM[28333] = 8'b0;
DRAM[28334] = 8'b100;
DRAM[28335] = 8'b111;
DRAM[28336] = 8'b0;
DRAM[28337] = 8'b11110;
DRAM[28338] = 8'b101101;
DRAM[28339] = 8'b1;
DRAM[28340] = 8'b100;
DRAM[28341] = 8'b111010;
DRAM[28342] = 8'b110101;
DRAM[28343] = 8'b10111;
DRAM[28344] = 8'b1010010;
DRAM[28345] = 8'b10000010;
DRAM[28346] = 8'b10100000;
DRAM[28347] = 8'b10010100;
DRAM[28348] = 8'b10001011;
DRAM[28349] = 8'b10011010;
DRAM[28350] = 8'b10100100;
DRAM[28351] = 8'b10011101;
DRAM[28352] = 8'b10010001;
DRAM[28353] = 8'b1111110;
DRAM[28354] = 8'b1111100;
DRAM[28355] = 8'b1101001;
DRAM[28356] = 8'b1010101;
DRAM[28357] = 8'b1001111;
DRAM[28358] = 8'b1000100;
DRAM[28359] = 8'b1000111;
DRAM[28360] = 8'b1000010;
DRAM[28361] = 8'b1100111;
DRAM[28362] = 8'b10001000;
DRAM[28363] = 8'b10010000;
DRAM[28364] = 8'b10100110;
DRAM[28365] = 8'b11000100;
DRAM[28366] = 8'b11010000;
DRAM[28367] = 8'b11011111;
DRAM[28368] = 8'b11111010;
DRAM[28369] = 8'b11111101;
DRAM[28370] = 8'b11110011;
DRAM[28371] = 8'b11110110;
DRAM[28372] = 8'b11100100;
DRAM[28373] = 8'b11011111;
DRAM[28374] = 8'b11010010;
DRAM[28375] = 8'b10110111;
DRAM[28376] = 8'b10101110;
DRAM[28377] = 8'b10011110;
DRAM[28378] = 8'b10011001;
DRAM[28379] = 8'b10010000;
DRAM[28380] = 8'b10001110;
DRAM[28381] = 8'b10011010;
DRAM[28382] = 8'b10010011;
DRAM[28383] = 8'b10011101;
DRAM[28384] = 8'b10011110;
DRAM[28385] = 8'b10111110;
DRAM[28386] = 8'b10111010;
DRAM[28387] = 8'b10001011;
DRAM[28388] = 8'b10101011;
DRAM[28389] = 8'b10000110;
DRAM[28390] = 8'b1111110;
DRAM[28391] = 8'b1111111;
DRAM[28392] = 8'b1111001;
DRAM[28393] = 8'b1110101;
DRAM[28394] = 8'b1110011;
DRAM[28395] = 8'b1110110;
DRAM[28396] = 8'b1110110;
DRAM[28397] = 8'b1110100;
DRAM[28398] = 8'b1110100;
DRAM[28399] = 8'b1110111;
DRAM[28400] = 8'b1110101;
DRAM[28401] = 8'b1110011;
DRAM[28402] = 8'b1110010;
DRAM[28403] = 8'b1110010;
DRAM[28404] = 8'b1110011;
DRAM[28405] = 8'b1110100;
DRAM[28406] = 8'b1110010;
DRAM[28407] = 8'b1110001;
DRAM[28408] = 8'b1110010;
DRAM[28409] = 8'b1110010;
DRAM[28410] = 8'b1110001;
DRAM[28411] = 8'b1110000;
DRAM[28412] = 8'b1101111;
DRAM[28413] = 8'b1101111;
DRAM[28414] = 8'b1101110;
DRAM[28415] = 8'b1101110;
DRAM[28416] = 8'b10000101;
DRAM[28417] = 8'b10000101;
DRAM[28418] = 8'b10000110;
DRAM[28419] = 8'b10000110;
DRAM[28420] = 8'b10000110;
DRAM[28421] = 8'b10000111;
DRAM[28422] = 8'b10000111;
DRAM[28423] = 8'b10000111;
DRAM[28424] = 8'b10000011;
DRAM[28425] = 8'b10000100;
DRAM[28426] = 8'b10000101;
DRAM[28427] = 8'b10000101;
DRAM[28428] = 8'b10000110;
DRAM[28429] = 8'b10000111;
DRAM[28430] = 8'b10001000;
DRAM[28431] = 8'b10001000;
DRAM[28432] = 8'b10001000;
DRAM[28433] = 8'b10001000;
DRAM[28434] = 8'b10001000;
DRAM[28435] = 8'b10001001;
DRAM[28436] = 8'b10001001;
DRAM[28437] = 8'b10001001;
DRAM[28438] = 8'b10001010;
DRAM[28439] = 8'b10001010;
DRAM[28440] = 8'b10001110;
DRAM[28441] = 8'b10001000;
DRAM[28442] = 8'b10001011;
DRAM[28443] = 8'b10010101;
DRAM[28444] = 8'b10010101;
DRAM[28445] = 8'b10001110;
DRAM[28446] = 8'b10010100;
DRAM[28447] = 8'b10100011;
DRAM[28448] = 8'b10010110;
DRAM[28449] = 8'b10100000;
DRAM[28450] = 8'b10111001;
DRAM[28451] = 8'b10110000;
DRAM[28452] = 8'b10111010;
DRAM[28453] = 8'b11010011;
DRAM[28454] = 8'b10111100;
DRAM[28455] = 8'b10101101;
DRAM[28456] = 8'b10100111;
DRAM[28457] = 8'b10101001;
DRAM[28458] = 8'b10001000;
DRAM[28459] = 8'b10011100;
DRAM[28460] = 8'b10010000;
DRAM[28461] = 8'b10010011;
DRAM[28462] = 8'b10011110;
DRAM[28463] = 8'b10100100;
DRAM[28464] = 8'b10011001;
DRAM[28465] = 8'b10110101;
DRAM[28466] = 8'b10100010;
DRAM[28467] = 8'b10011110;
DRAM[28468] = 8'b10011001;
DRAM[28469] = 8'b10100011;
DRAM[28470] = 8'b10100000;
DRAM[28471] = 8'b11000101;
DRAM[28472] = 8'b11001110;
DRAM[28473] = 8'b10111000;
DRAM[28474] = 8'b11011001;
DRAM[28475] = 8'b11100001;
DRAM[28476] = 8'b11001001;
DRAM[28477] = 8'b11101111;
DRAM[28478] = 8'b11011000;
DRAM[28479] = 8'b11011000;
DRAM[28480] = 8'b11101001;
DRAM[28481] = 8'b11011101;
DRAM[28482] = 8'b11000000;
DRAM[28483] = 8'b11010111;
DRAM[28484] = 8'b10111101;
DRAM[28485] = 8'b10111100;
DRAM[28486] = 8'b10111001;
DRAM[28487] = 8'b10011110;
DRAM[28488] = 8'b10010100;
DRAM[28489] = 8'b1100000;
DRAM[28490] = 8'b1010001;
DRAM[28491] = 8'b1010001;
DRAM[28492] = 8'b1100110;
DRAM[28493] = 8'b1100001;
DRAM[28494] = 8'b1111010;
DRAM[28495] = 8'b10000001;
DRAM[28496] = 8'b10010000;
DRAM[28497] = 8'b10100110;
DRAM[28498] = 8'b10110010;
DRAM[28499] = 8'b10110100;
DRAM[28500] = 8'b10110110;
DRAM[28501] = 8'b10110110;
DRAM[28502] = 8'b11000000;
DRAM[28503] = 8'b11010100;
DRAM[28504] = 8'b11011001;
DRAM[28505] = 8'b11001011;
DRAM[28506] = 8'b11001101;
DRAM[28507] = 8'b11011101;
DRAM[28508] = 8'b11011100;
DRAM[28509] = 8'b11001000;
DRAM[28510] = 8'b10111111;
DRAM[28511] = 8'b11000110;
DRAM[28512] = 8'b10111111;
DRAM[28513] = 8'b11001111;
DRAM[28514] = 8'b11000111;
DRAM[28515] = 8'b10100011;
DRAM[28516] = 8'b10001010;
DRAM[28517] = 8'b10000101;
DRAM[28518] = 8'b1111000;
DRAM[28519] = 8'b1100010;
DRAM[28520] = 8'b1100001;
DRAM[28521] = 8'b1101100;
DRAM[28522] = 8'b10001000;
DRAM[28523] = 8'b1110100;
DRAM[28524] = 8'b1100111;
DRAM[28525] = 8'b1100101;
DRAM[28526] = 8'b111110;
DRAM[28527] = 8'b101110;
DRAM[28528] = 8'b110100;
DRAM[28529] = 8'b111000;
DRAM[28530] = 8'b111111;
DRAM[28531] = 8'b1010001;
DRAM[28532] = 8'b1100000;
DRAM[28533] = 8'b1011100;
DRAM[28534] = 8'b1011000;
DRAM[28535] = 8'b1100010;
DRAM[28536] = 8'b1101000;
DRAM[28537] = 8'b1100010;
DRAM[28538] = 8'b1111000;
DRAM[28539] = 8'b1111100;
DRAM[28540] = 8'b10000100;
DRAM[28541] = 8'b1111100;
DRAM[28542] = 8'b10001101;
DRAM[28543] = 8'b10001101;
DRAM[28544] = 8'b10010111;
DRAM[28545] = 8'b10001010;
DRAM[28546] = 8'b10010010;
DRAM[28547] = 8'b10011110;
DRAM[28548] = 8'b10001100;
DRAM[28549] = 8'b10010011;
DRAM[28550] = 8'b10110011;
DRAM[28551] = 8'b10110000;
DRAM[28552] = 8'b10111000;
DRAM[28553] = 8'b10101011;
DRAM[28554] = 8'b10110001;
DRAM[28555] = 8'b10111001;
DRAM[28556] = 8'b10110110;
DRAM[28557] = 8'b10111111;
DRAM[28558] = 8'b11000010;
DRAM[28559] = 8'b10110000;
DRAM[28560] = 8'b10111101;
DRAM[28561] = 8'b10101101;
DRAM[28562] = 8'b10101110;
DRAM[28563] = 8'b11000001;
DRAM[28564] = 8'b10011110;
DRAM[28565] = 8'b10100111;
DRAM[28566] = 8'b10101001;
DRAM[28567] = 8'b10100100;
DRAM[28568] = 8'b10100000;
DRAM[28569] = 8'b10011101;
DRAM[28570] = 8'b10100100;
DRAM[28571] = 8'b10011111;
DRAM[28572] = 8'b10010000;
DRAM[28573] = 8'b10010001;
DRAM[28574] = 8'b10000111;
DRAM[28575] = 8'b1100101;
DRAM[28576] = 8'b1010101;
DRAM[28577] = 8'b1000001;
DRAM[28578] = 8'b100111;
DRAM[28579] = 8'b10110;
DRAM[28580] = 8'b10100;
DRAM[28581] = 8'b10110;
DRAM[28582] = 8'b10001;
DRAM[28583] = 8'b111;
DRAM[28584] = 8'b10011;
DRAM[28585] = 8'b1010;
DRAM[28586] = 8'b100;
DRAM[28587] = 8'b1100;
DRAM[28588] = 8'b1001;
DRAM[28589] = 8'b1;
DRAM[28590] = 8'b1010;
DRAM[28591] = 8'b1;
DRAM[28592] = 8'b100;
DRAM[28593] = 8'b10000;
DRAM[28594] = 8'b100101;
DRAM[28595] = 8'b10001;
DRAM[28596] = 8'b1000;
DRAM[28597] = 8'b10001;
DRAM[28598] = 8'b10101;
DRAM[28599] = 8'b111010;
DRAM[28600] = 8'b1110010;
DRAM[28601] = 8'b10000111;
DRAM[28602] = 8'b10011110;
DRAM[28603] = 8'b10100111;
DRAM[28604] = 8'b10100001;
DRAM[28605] = 8'b10011000;
DRAM[28606] = 8'b10010010;
DRAM[28607] = 8'b10010001;
DRAM[28608] = 8'b10001111;
DRAM[28609] = 8'b1111100;
DRAM[28610] = 8'b1111101;
DRAM[28611] = 8'b1101010;
DRAM[28612] = 8'b1010100;
DRAM[28613] = 8'b1010000;
DRAM[28614] = 8'b1001000;
DRAM[28615] = 8'b1001001;
DRAM[28616] = 8'b1001111;
DRAM[28617] = 8'b1010000;
DRAM[28618] = 8'b10000010;
DRAM[28619] = 8'b10001111;
DRAM[28620] = 8'b10100010;
DRAM[28621] = 8'b10111000;
DRAM[28622] = 8'b10110101;
DRAM[28623] = 8'b11101001;
DRAM[28624] = 8'b11101111;
DRAM[28625] = 8'b11110110;
DRAM[28626] = 8'b11110000;
DRAM[28627] = 8'b11111111;
DRAM[28628] = 8'b11110010;
DRAM[28629] = 8'b11011000;
DRAM[28630] = 8'b11011010;
DRAM[28631] = 8'b11000011;
DRAM[28632] = 8'b10101110;
DRAM[28633] = 8'b10010100;
DRAM[28634] = 8'b10011011;
DRAM[28635] = 8'b10001010;
DRAM[28636] = 8'b10010111;
DRAM[28637] = 8'b10010000;
DRAM[28638] = 8'b10010111;
DRAM[28639] = 8'b10100011;
DRAM[28640] = 8'b10011111;
DRAM[28641] = 8'b11000010;
DRAM[28642] = 8'b10111100;
DRAM[28643] = 8'b1111000;
DRAM[28644] = 8'b10100010;
DRAM[28645] = 8'b10000101;
DRAM[28646] = 8'b1110001;
DRAM[28647] = 8'b1111101;
DRAM[28648] = 8'b10000001;
DRAM[28649] = 8'b1111011;
DRAM[28650] = 8'b1111000;
DRAM[28651] = 8'b1111001;
DRAM[28652] = 8'b1110111;
DRAM[28653] = 8'b1110100;
DRAM[28654] = 8'b1110011;
DRAM[28655] = 8'b1110110;
DRAM[28656] = 8'b1110101;
DRAM[28657] = 8'b1110100;
DRAM[28658] = 8'b1110010;
DRAM[28659] = 8'b1110010;
DRAM[28660] = 8'b1110100;
DRAM[28661] = 8'b1110100;
DRAM[28662] = 8'b1110010;
DRAM[28663] = 8'b1110001;
DRAM[28664] = 8'b1110010;
DRAM[28665] = 8'b1110010;
DRAM[28666] = 8'b1110001;
DRAM[28667] = 8'b1110000;
DRAM[28668] = 8'b1110000;
DRAM[28669] = 8'b1101111;
DRAM[28670] = 8'b1101110;
DRAM[28671] = 8'b1101110;
DRAM[28672] = 8'b10000100;
DRAM[28673] = 8'b10000100;
DRAM[28674] = 8'b10000100;
DRAM[28675] = 8'b10000101;
DRAM[28676] = 8'b10000101;
DRAM[28677] = 8'b10000101;
DRAM[28678] = 8'b10000110;
DRAM[28679] = 8'b10000110;
DRAM[28680] = 8'b10001000;
DRAM[28681] = 8'b10001000;
DRAM[28682] = 8'b10001000;
DRAM[28683] = 8'b10001001;
DRAM[28684] = 8'b10001001;
DRAM[28685] = 8'b10001010;
DRAM[28686] = 8'b10001010;
DRAM[28687] = 8'b10001010;
DRAM[28688] = 8'b10001011;
DRAM[28689] = 8'b10001010;
DRAM[28690] = 8'b10001010;
DRAM[28691] = 8'b10001001;
DRAM[28692] = 8'b10001001;
DRAM[28693] = 8'b10001010;
DRAM[28694] = 8'b10001010;
DRAM[28695] = 8'b10001011;
DRAM[28696] = 8'b10001100;
DRAM[28697] = 8'b10001100;
DRAM[28698] = 8'b10001101;
DRAM[28699] = 8'b10001110;
DRAM[28700] = 8'b10001110;
DRAM[28701] = 8'b10001111;
DRAM[28702] = 8'b10010000;
DRAM[28703] = 8'b10010000;
DRAM[28704] = 8'b10010110;
DRAM[28705] = 8'b10011111;
DRAM[28706] = 8'b10011100;
DRAM[28707] = 8'b10100010;
DRAM[28708] = 8'b10111100;
DRAM[28709] = 8'b11001010;
DRAM[28710] = 8'b10111111;
DRAM[28711] = 8'b10110010;
DRAM[28712] = 8'b10110000;
DRAM[28713] = 8'b10011010;
DRAM[28714] = 8'b10100110;
DRAM[28715] = 8'b10100100;
DRAM[28716] = 8'b10010011;
DRAM[28717] = 8'b10010111;
DRAM[28718] = 8'b10011000;
DRAM[28719] = 8'b10011010;
DRAM[28720] = 8'b10100000;
DRAM[28721] = 8'b10011110;
DRAM[28722] = 8'b10011111;
DRAM[28723] = 8'b10100010;
DRAM[28724] = 8'b10100000;
DRAM[28725] = 8'b10100000;
DRAM[28726] = 8'b10101101;
DRAM[28727] = 8'b10111111;
DRAM[28728] = 8'b11000101;
DRAM[28729] = 8'b11000001;
DRAM[28730] = 8'b11011011;
DRAM[28731] = 8'b11010001;
DRAM[28732] = 8'b11100110;
DRAM[28733] = 8'b11100111;
DRAM[28734] = 8'b11100100;
DRAM[28735] = 8'b11011110;
DRAM[28736] = 8'b11101110;
DRAM[28737] = 8'b11011110;
DRAM[28738] = 8'b10111011;
DRAM[28739] = 8'b11100001;
DRAM[28740] = 8'b10110101;
DRAM[28741] = 8'b10111010;
DRAM[28742] = 8'b10110111;
DRAM[28743] = 8'b10100001;
DRAM[28744] = 8'b10000011;
DRAM[28745] = 8'b1100001;
DRAM[28746] = 8'b1001111;
DRAM[28747] = 8'b1011110;
DRAM[28748] = 8'b1101101;
DRAM[28749] = 8'b1101101;
DRAM[28750] = 8'b1110000;
DRAM[28751] = 8'b1111011;
DRAM[28752] = 8'b10001011;
DRAM[28753] = 8'b10100101;
DRAM[28754] = 8'b10110000;
DRAM[28755] = 8'b10101110;
DRAM[28756] = 8'b10110111;
DRAM[28757] = 8'b11000011;
DRAM[28758] = 8'b11001011;
DRAM[28759] = 8'b11010100;
DRAM[28760] = 8'b11001011;
DRAM[28761] = 8'b11000110;
DRAM[28762] = 8'b11010111;
DRAM[28763] = 8'b11011100;
DRAM[28764] = 8'b11001100;
DRAM[28765] = 8'b11010001;
DRAM[28766] = 8'b11010000;
DRAM[28767] = 8'b10110000;
DRAM[28768] = 8'b10101100;
DRAM[28769] = 8'b10110100;
DRAM[28770] = 8'b10100011;
DRAM[28771] = 8'b10010011;
DRAM[28772] = 8'b1111001;
DRAM[28773] = 8'b10000011;
DRAM[28774] = 8'b1111100;
DRAM[28775] = 8'b10011010;
DRAM[28776] = 8'b11000110;
DRAM[28777] = 8'b10011001;
DRAM[28778] = 8'b10011001;
DRAM[28779] = 8'b1111000;
DRAM[28780] = 8'b1010011;
DRAM[28781] = 8'b1001110;
DRAM[28782] = 8'b101111;
DRAM[28783] = 8'b101011;
DRAM[28784] = 8'b101101;
DRAM[28785] = 8'b11101;
DRAM[28786] = 8'b110001;
DRAM[28787] = 8'b1001000;
DRAM[28788] = 8'b1000101;
DRAM[28789] = 8'b1010010;
DRAM[28790] = 8'b1011111;
DRAM[28791] = 8'b1001111;
DRAM[28792] = 8'b1011100;
DRAM[28793] = 8'b1101000;
DRAM[28794] = 8'b1110001;
DRAM[28795] = 8'b1110010;
DRAM[28796] = 8'b1110110;
DRAM[28797] = 8'b10000001;
DRAM[28798] = 8'b10001100;
DRAM[28799] = 8'b10001111;
DRAM[28800] = 8'b10011000;
DRAM[28801] = 8'b10100000;
DRAM[28802] = 8'b10011010;
DRAM[28803] = 8'b10010100;
DRAM[28804] = 8'b10011100;
DRAM[28805] = 8'b10100011;
DRAM[28806] = 8'b10101000;
DRAM[28807] = 8'b10110001;
DRAM[28808] = 8'b10111010;
DRAM[28809] = 8'b10101110;
DRAM[28810] = 8'b11001010;
DRAM[28811] = 8'b10111011;
DRAM[28812] = 8'b10111110;
DRAM[28813] = 8'b10110110;
DRAM[28814] = 8'b10111110;
DRAM[28815] = 8'b10111110;
DRAM[28816] = 8'b11001011;
DRAM[28817] = 8'b10111110;
DRAM[28818] = 8'b10110000;
DRAM[28819] = 8'b10100111;
DRAM[28820] = 8'b10100111;
DRAM[28821] = 8'b10101001;
DRAM[28822] = 8'b10101001;
DRAM[28823] = 8'b10100111;
DRAM[28824] = 8'b10010010;
DRAM[28825] = 8'b10011000;
DRAM[28826] = 8'b10101101;
DRAM[28827] = 8'b10010111;
DRAM[28828] = 8'b10011100;
DRAM[28829] = 8'b10100001;
DRAM[28830] = 8'b10100001;
DRAM[28831] = 8'b1101100;
DRAM[28832] = 8'b1010000;
DRAM[28833] = 8'b1001101;
DRAM[28834] = 8'b101010;
DRAM[28835] = 8'b111000;
DRAM[28836] = 8'b11011;
DRAM[28837] = 8'b10001;
DRAM[28838] = 8'b10001;
DRAM[28839] = 8'b1;
DRAM[28840] = 8'b1110;
DRAM[28841] = 8'b1101;
DRAM[28842] = 8'b1001;
DRAM[28843] = 8'b100;
DRAM[28844] = 8'b10;
DRAM[28845] = 8'b11;
DRAM[28846] = 8'b11;
DRAM[28847] = 8'b10;
DRAM[28848] = 8'b1000;
DRAM[28849] = 8'b1110;
DRAM[28850] = 8'b10101;
DRAM[28851] = 8'b1100;
DRAM[28852] = 8'b11100;
DRAM[28853] = 8'b110010;
DRAM[28854] = 8'b110001;
DRAM[28855] = 8'b111100;
DRAM[28856] = 8'b1101101;
DRAM[28857] = 8'b10010110;
DRAM[28858] = 8'b10101010;
DRAM[28859] = 8'b10011111;
DRAM[28860] = 8'b10010011;
DRAM[28861] = 8'b10001101;
DRAM[28862] = 8'b10001011;
DRAM[28863] = 8'b10001111;
DRAM[28864] = 8'b10001101;
DRAM[28865] = 8'b10000100;
DRAM[28866] = 8'b1110111;
DRAM[28867] = 8'b1101010;
DRAM[28868] = 8'b1100000;
DRAM[28869] = 8'b1011000;
DRAM[28870] = 8'b1010010;
DRAM[28871] = 8'b1001110;
DRAM[28872] = 8'b1011011;
DRAM[28873] = 8'b1010101;
DRAM[28874] = 8'b1101111;
DRAM[28875] = 8'b10011001;
DRAM[28876] = 8'b1110111;
DRAM[28877] = 8'b10101010;
DRAM[28878] = 8'b11011011;
DRAM[28879] = 8'b11000000;
DRAM[28880] = 8'b11101100;
DRAM[28881] = 8'b11110000;
DRAM[28882] = 8'b11111011;
DRAM[28883] = 8'b11101110;
DRAM[28884] = 8'b11110111;
DRAM[28885] = 8'b11100110;
DRAM[28886] = 8'b11010110;
DRAM[28887] = 8'b10111000;
DRAM[28888] = 8'b10110101;
DRAM[28889] = 8'b10011001;
DRAM[28890] = 8'b10011101;
DRAM[28891] = 8'b10010011;
DRAM[28892] = 8'b10001111;
DRAM[28893] = 8'b10010111;
DRAM[28894] = 8'b10010110;
DRAM[28895] = 8'b10110111;
DRAM[28896] = 8'b10111010;
DRAM[28897] = 8'b10101000;
DRAM[28898] = 8'b10100001;
DRAM[28899] = 8'b10010010;
DRAM[28900] = 8'b10001110;
DRAM[28901] = 8'b10001101;
DRAM[28902] = 8'b1111001;
DRAM[28903] = 8'b1110101;
DRAM[28904] = 8'b1110111;
DRAM[28905] = 8'b1111000;
DRAM[28906] = 8'b1111001;
DRAM[28907] = 8'b1111010;
DRAM[28908] = 8'b1111001;
DRAM[28909] = 8'b1111000;
DRAM[28910] = 8'b1110111;
DRAM[28911] = 8'b1110110;
DRAM[28912] = 8'b1110101;
DRAM[28913] = 8'b1110100;
DRAM[28914] = 8'b1110011;
DRAM[28915] = 8'b1110100;
DRAM[28916] = 8'b1110101;
DRAM[28917] = 8'b1110101;
DRAM[28918] = 8'b1110011;
DRAM[28919] = 8'b1110001;
DRAM[28920] = 8'b1110011;
DRAM[28921] = 8'b1110011;
DRAM[28922] = 8'b1110011;
DRAM[28923] = 8'b1110010;
DRAM[28924] = 8'b1110010;
DRAM[28925] = 8'b1110001;
DRAM[28926] = 8'b1110001;
DRAM[28927] = 8'b1110001;
DRAM[28928] = 8'b10000100;
DRAM[28929] = 8'b10000100;
DRAM[28930] = 8'b10000101;
DRAM[28931] = 8'b10000101;
DRAM[28932] = 8'b10000101;
DRAM[28933] = 8'b10000110;
DRAM[28934] = 8'b10000110;
DRAM[28935] = 8'b10000110;
DRAM[28936] = 8'b10001000;
DRAM[28937] = 8'b10001000;
DRAM[28938] = 8'b10001001;
DRAM[28939] = 8'b10001001;
DRAM[28940] = 8'b10001001;
DRAM[28941] = 8'b10001010;
DRAM[28942] = 8'b10001010;
DRAM[28943] = 8'b10001010;
DRAM[28944] = 8'b10001011;
DRAM[28945] = 8'b10001010;
DRAM[28946] = 8'b10001010;
DRAM[28947] = 8'b10001001;
DRAM[28948] = 8'b10001001;
DRAM[28949] = 8'b10001010;
DRAM[28950] = 8'b10001010;
DRAM[28951] = 8'b10001011;
DRAM[28952] = 8'b10001100;
DRAM[28953] = 8'b10001100;
DRAM[28954] = 8'b10001101;
DRAM[28955] = 8'b10001110;
DRAM[28956] = 8'b10001110;
DRAM[28957] = 8'b10001111;
DRAM[28958] = 8'b10010000;
DRAM[28959] = 8'b10010000;
DRAM[28960] = 8'b10010011;
DRAM[28961] = 8'b10010110;
DRAM[28962] = 8'b10011000;
DRAM[28963] = 8'b10101001;
DRAM[28964] = 8'b11000011;
DRAM[28965] = 8'b11001000;
DRAM[28966] = 8'b11000000;
DRAM[28967] = 8'b11000000;
DRAM[28968] = 8'b10110010;
DRAM[28969] = 8'b10100100;
DRAM[28970] = 8'b10101101;
DRAM[28971] = 8'b10100101;
DRAM[28972] = 8'b10011000;
DRAM[28973] = 8'b10011010;
DRAM[28974] = 8'b10011010;
DRAM[28975] = 8'b10100101;
DRAM[28976] = 8'b10010110;
DRAM[28977] = 8'b10010101;
DRAM[28978] = 8'b10011001;
DRAM[28979] = 8'b10011110;
DRAM[28980] = 8'b10011110;
DRAM[28981] = 8'b10011110;
DRAM[28982] = 8'b10101100;
DRAM[28983] = 8'b10111101;
DRAM[28984] = 8'b11000100;
DRAM[28985] = 8'b11000110;
DRAM[28986] = 8'b11011100;
DRAM[28987] = 8'b11010111;
DRAM[28988] = 8'b11100001;
DRAM[28989] = 8'b11100111;
DRAM[28990] = 8'b11100001;
DRAM[28991] = 8'b11100001;
DRAM[28992] = 8'b11110010;
DRAM[28993] = 8'b11011010;
DRAM[28994] = 8'b11010100;
DRAM[28995] = 8'b11010011;
DRAM[28996] = 8'b10111100;
DRAM[28997] = 8'b10110000;
DRAM[28998] = 8'b10111001;
DRAM[28999] = 8'b10011101;
DRAM[29000] = 8'b1110111;
DRAM[29001] = 8'b1011010;
DRAM[29002] = 8'b1001010;
DRAM[29003] = 8'b1010110;
DRAM[29004] = 8'b1100011;
DRAM[29005] = 8'b1100110;
DRAM[29006] = 8'b1110000;
DRAM[29007] = 8'b10000000;
DRAM[29008] = 8'b10001001;
DRAM[29009] = 8'b10011110;
DRAM[29010] = 8'b10100111;
DRAM[29011] = 8'b10100111;
DRAM[29012] = 8'b10110010;
DRAM[29013] = 8'b10111011;
DRAM[29014] = 8'b10111101;
DRAM[29015] = 8'b11000000;
DRAM[29016] = 8'b11010101;
DRAM[29017] = 8'b11011001;
DRAM[29018] = 8'b11001101;
DRAM[29019] = 8'b11001111;
DRAM[29020] = 8'b11011011;
DRAM[29021] = 8'b10111111;
DRAM[29022] = 8'b10100001;
DRAM[29023] = 8'b10101100;
DRAM[29024] = 8'b11000011;
DRAM[29025] = 8'b10111111;
DRAM[29026] = 8'b10001010;
DRAM[29027] = 8'b10001001;
DRAM[29028] = 8'b10100100;
DRAM[29029] = 8'b11000011;
DRAM[29030] = 8'b10111001;
DRAM[29031] = 8'b11000011;
DRAM[29032] = 8'b10110010;
DRAM[29033] = 8'b1101101;
DRAM[29034] = 8'b1010001;
DRAM[29035] = 8'b101011;
DRAM[29036] = 8'b101011;
DRAM[29037] = 8'b10111;
DRAM[29038] = 8'b10000;
DRAM[29039] = 8'b1101;
DRAM[29040] = 8'b11000;
DRAM[29041] = 8'b1100;
DRAM[29042] = 8'b100010;
DRAM[29043] = 8'b1000110;
DRAM[29044] = 8'b1010000;
DRAM[29045] = 8'b1010000;
DRAM[29046] = 8'b1010001;
DRAM[29047] = 8'b1001011;
DRAM[29048] = 8'b1010110;
DRAM[29049] = 8'b1011111;
DRAM[29050] = 8'b1101011;
DRAM[29051] = 8'b1110101;
DRAM[29052] = 8'b1111111;
DRAM[29053] = 8'b10001001;
DRAM[29054] = 8'b10001111;
DRAM[29055] = 8'b10010000;
DRAM[29056] = 8'b10010010;
DRAM[29057] = 8'b10011011;
DRAM[29058] = 8'b10011000;
DRAM[29059] = 8'b10010101;
DRAM[29060] = 8'b10011111;
DRAM[29061] = 8'b10101000;
DRAM[29062] = 8'b10101101;
DRAM[29063] = 8'b10110110;
DRAM[29064] = 8'b10111110;
DRAM[29065] = 8'b10101110;
DRAM[29066] = 8'b11000101;
DRAM[29067] = 8'b10111010;
DRAM[29068] = 8'b11000001;
DRAM[29069] = 8'b10111101;
DRAM[29070] = 8'b10111101;
DRAM[29071] = 8'b10111000;
DRAM[29072] = 8'b10111111;
DRAM[29073] = 8'b10111100;
DRAM[29074] = 8'b10110111;
DRAM[29075] = 8'b10110010;
DRAM[29076] = 8'b10101101;
DRAM[29077] = 8'b10101001;
DRAM[29078] = 8'b10100101;
DRAM[29079] = 8'b10100010;
DRAM[29080] = 8'b10011011;
DRAM[29081] = 8'b10011111;
DRAM[29082] = 8'b10100101;
DRAM[29083] = 8'b10100101;
DRAM[29084] = 8'b10001111;
DRAM[29085] = 8'b10100110;
DRAM[29086] = 8'b10010000;
DRAM[29087] = 8'b10001100;
DRAM[29088] = 8'b1101111;
DRAM[29089] = 8'b1010111;
DRAM[29090] = 8'b1000100;
DRAM[29091] = 8'b111100;
DRAM[29092] = 8'b100110;
DRAM[29093] = 8'b100000;
DRAM[29094] = 8'b1111;
DRAM[29095] = 8'b1100;
DRAM[29096] = 8'b10100;
DRAM[29097] = 8'b10010;
DRAM[29098] = 8'b1111;
DRAM[29099] = 8'b1011;
DRAM[29100] = 8'b1001;
DRAM[29101] = 8'b1001;
DRAM[29102] = 8'b1001;
DRAM[29103] = 8'b1000;
DRAM[29104] = 8'b1010;
DRAM[29105] = 8'b1010;
DRAM[29106] = 8'b10010;
DRAM[29107] = 8'b1101;
DRAM[29108] = 8'b10100;
DRAM[29109] = 8'b100011;
DRAM[29110] = 8'b110111;
DRAM[29111] = 8'b1100011;
DRAM[29112] = 8'b10000100;
DRAM[29113] = 8'b10100100;
DRAM[29114] = 8'b10110001;
DRAM[29115] = 8'b10101000;
DRAM[29116] = 8'b10100010;
DRAM[29117] = 8'b10011011;
DRAM[29118] = 8'b10001111;
DRAM[29119] = 8'b10001010;
DRAM[29120] = 8'b10000010;
DRAM[29121] = 8'b1111100;
DRAM[29122] = 8'b1110010;
DRAM[29123] = 8'b1100111;
DRAM[29124] = 8'b1011110;
DRAM[29125] = 8'b1010111;
DRAM[29126] = 8'b1010011;
DRAM[29127] = 8'b1010001;
DRAM[29128] = 8'b1011000;
DRAM[29129] = 8'b1100000;
DRAM[29130] = 8'b1100000;
DRAM[29131] = 8'b10000110;
DRAM[29132] = 8'b10001010;
DRAM[29133] = 8'b10011001;
DRAM[29134] = 8'b11001011;
DRAM[29135] = 8'b11001010;
DRAM[29136] = 8'b11100101;
DRAM[29137] = 8'b11101100;
DRAM[29138] = 8'b11111011;
DRAM[29139] = 8'b11110001;
DRAM[29140] = 8'b11111010;
DRAM[29141] = 8'b11101000;
DRAM[29142] = 8'b11011000;
DRAM[29143] = 8'b10111100;
DRAM[29144] = 8'b10111000;
DRAM[29145] = 8'b10011101;
DRAM[29146] = 8'b10010010;
DRAM[29147] = 8'b10011011;
DRAM[29148] = 8'b10011000;
DRAM[29149] = 8'b10011101;
DRAM[29150] = 8'b10011110;
DRAM[29151] = 8'b10111011;
DRAM[29152] = 8'b10111101;
DRAM[29153] = 8'b10100110;
DRAM[29154] = 8'b10011001;
DRAM[29155] = 8'b10000101;
DRAM[29156] = 8'b10000010;
DRAM[29157] = 8'b10001000;
DRAM[29158] = 8'b1111100;
DRAM[29159] = 8'b1111110;
DRAM[29160] = 8'b1111000;
DRAM[29161] = 8'b1111000;
DRAM[29162] = 8'b1111001;
DRAM[29163] = 8'b1111010;
DRAM[29164] = 8'b1111001;
DRAM[29165] = 8'b1111000;
DRAM[29166] = 8'b1110111;
DRAM[29167] = 8'b1110110;
DRAM[29168] = 8'b1110110;
DRAM[29169] = 8'b1110101;
DRAM[29170] = 8'b1110100;
DRAM[29171] = 8'b1110100;
DRAM[29172] = 8'b1110110;
DRAM[29173] = 8'b1110101;
DRAM[29174] = 8'b1110011;
DRAM[29175] = 8'b1110001;
DRAM[29176] = 8'b1110011;
DRAM[29177] = 8'b1110011;
DRAM[29178] = 8'b1110011;
DRAM[29179] = 8'b1110010;
DRAM[29180] = 8'b1110010;
DRAM[29181] = 8'b1110010;
DRAM[29182] = 8'b1110001;
DRAM[29183] = 8'b1110001;
DRAM[29184] = 8'b10000101;
DRAM[29185] = 8'b10000101;
DRAM[29186] = 8'b10000101;
DRAM[29187] = 8'b10000110;
DRAM[29188] = 8'b10000110;
DRAM[29189] = 8'b10000110;
DRAM[29190] = 8'b10000111;
DRAM[29191] = 8'b10000111;
DRAM[29192] = 8'b10001000;
DRAM[29193] = 8'b10001001;
DRAM[29194] = 8'b10001001;
DRAM[29195] = 8'b10001001;
DRAM[29196] = 8'b10001010;
DRAM[29197] = 8'b10001010;
DRAM[29198] = 8'b10001010;
DRAM[29199] = 8'b10001010;
DRAM[29200] = 8'b10001011;
DRAM[29201] = 8'b10001011;
DRAM[29202] = 8'b10001010;
DRAM[29203] = 8'b10001010;
DRAM[29204] = 8'b10001010;
DRAM[29205] = 8'b10001010;
DRAM[29206] = 8'b10001011;
DRAM[29207] = 8'b10001011;
DRAM[29208] = 8'b10001100;
DRAM[29209] = 8'b10001100;
DRAM[29210] = 8'b10001101;
DRAM[29211] = 8'b10001110;
DRAM[29212] = 8'b10001110;
DRAM[29213] = 8'b10001111;
DRAM[29214] = 8'b10010000;
DRAM[29215] = 8'b10010000;
DRAM[29216] = 8'b10010001;
DRAM[29217] = 8'b10010001;
DRAM[29218] = 8'b10010111;
DRAM[29219] = 8'b10101101;
DRAM[29220] = 8'b11000100;
DRAM[29221] = 8'b11000001;
DRAM[29222] = 8'b10111101;
DRAM[29223] = 8'b11000111;
DRAM[29224] = 8'b10110010;
DRAM[29225] = 8'b10101101;
DRAM[29226] = 8'b10101101;
DRAM[29227] = 8'b10011101;
DRAM[29228] = 8'b10010111;
DRAM[29229] = 8'b10010111;
DRAM[29230] = 8'b10010010;
DRAM[29231] = 8'b10100111;
DRAM[29232] = 8'b10001100;
DRAM[29233] = 8'b10001101;
DRAM[29234] = 8'b10010100;
DRAM[29235] = 8'b10011101;
DRAM[29236] = 8'b10011111;
DRAM[29237] = 8'b10100000;
DRAM[29238] = 8'b10101110;
DRAM[29239] = 8'b10111111;
DRAM[29240] = 8'b11000010;
DRAM[29241] = 8'b11001010;
DRAM[29242] = 8'b11011010;
DRAM[29243] = 8'b11011110;
DRAM[29244] = 8'b11011011;
DRAM[29245] = 8'b11101001;
DRAM[29246] = 8'b11011101;
DRAM[29247] = 8'b11100011;
DRAM[29248] = 8'b11110001;
DRAM[29249] = 8'b11011010;
DRAM[29250] = 8'b11100001;
DRAM[29251] = 8'b11001101;
DRAM[29252] = 8'b10110001;
DRAM[29253] = 8'b10110011;
DRAM[29254] = 8'b10110000;
DRAM[29255] = 8'b10010101;
DRAM[29256] = 8'b1100101;
DRAM[29257] = 8'b1010011;
DRAM[29258] = 8'b1001100;
DRAM[29259] = 8'b1010111;
DRAM[29260] = 8'b1100000;
DRAM[29261] = 8'b1100011;
DRAM[29262] = 8'b1110000;
DRAM[29263] = 8'b10000011;
DRAM[29264] = 8'b10001110;
DRAM[29265] = 8'b10100001;
DRAM[29266] = 8'b10101000;
DRAM[29267] = 8'b10101011;
DRAM[29268] = 8'b10110111;
DRAM[29269] = 8'b10111011;
DRAM[29270] = 8'b10110101;
DRAM[29271] = 8'b10110011;
DRAM[29272] = 8'b10110000;
DRAM[29273] = 8'b11000100;
DRAM[29274] = 8'b11000111;
DRAM[29275] = 8'b11001011;
DRAM[29276] = 8'b11010001;
DRAM[29277] = 8'b10110100;
DRAM[29278] = 8'b10011110;
DRAM[29279] = 8'b10110001;
DRAM[29280] = 8'b10000101;
DRAM[29281] = 8'b1111110;
DRAM[29282] = 8'b10001111;
DRAM[29283] = 8'b11001111;
DRAM[29284] = 8'b11000010;
DRAM[29285] = 8'b10110001;
DRAM[29286] = 8'b10100100;
DRAM[29287] = 8'b1110000;
DRAM[29288] = 8'b111011;
DRAM[29289] = 8'b110010;
DRAM[29290] = 8'b1110;
DRAM[29291] = 8'b11;
DRAM[29292] = 8'b0;
DRAM[29293] = 8'b0;
DRAM[29294] = 8'b0;
DRAM[29295] = 8'b0;
DRAM[29296] = 8'b10;
DRAM[29297] = 8'b0;
DRAM[29298] = 8'b1101;
DRAM[29299] = 8'b110010;
DRAM[29300] = 8'b1001101;
DRAM[29301] = 8'b1001000;
DRAM[29302] = 8'b1000001;
DRAM[29303] = 8'b1001010;
DRAM[29304] = 8'b1010000;
DRAM[29305] = 8'b1010101;
DRAM[29306] = 8'b1100100;
DRAM[29307] = 8'b1111001;
DRAM[29308] = 8'b10001010;
DRAM[29309] = 8'b10010001;
DRAM[29310] = 8'b10010011;
DRAM[29311] = 8'b10010011;
DRAM[29312] = 8'b10010010;
DRAM[29313] = 8'b10011101;
DRAM[29314] = 8'b10011100;
DRAM[29315] = 8'b10011011;
DRAM[29316] = 8'b10100111;
DRAM[29317] = 8'b10101111;
DRAM[29318] = 8'b10110011;
DRAM[29319] = 8'b10111100;
DRAM[29320] = 8'b11000100;
DRAM[29321] = 8'b10110010;
DRAM[29322] = 8'b11000010;
DRAM[29323] = 8'b10111011;
DRAM[29324] = 8'b11000100;
DRAM[29325] = 8'b11000111;
DRAM[29326] = 8'b11000001;
DRAM[29327] = 8'b10110111;
DRAM[29328] = 8'b10111001;
DRAM[29329] = 8'b10111011;
DRAM[29330] = 8'b10111100;
DRAM[29331] = 8'b10111000;
DRAM[29332] = 8'b10110010;
DRAM[29333] = 8'b10101100;
DRAM[29334] = 8'b10101001;
DRAM[29335] = 8'b10101001;
DRAM[29336] = 8'b10100000;
DRAM[29337] = 8'b10100001;
DRAM[29338] = 8'b10100011;
DRAM[29339] = 8'b10100110;
DRAM[29340] = 8'b10010011;
DRAM[29341] = 8'b10011101;
DRAM[29342] = 8'b10001010;
DRAM[29343] = 8'b10101011;
DRAM[29344] = 8'b10001001;
DRAM[29345] = 8'b1011100;
DRAM[29346] = 8'b1010111;
DRAM[29347] = 8'b111001;
DRAM[29348] = 8'b110011;
DRAM[29349] = 8'b101001;
DRAM[29350] = 8'b1110;
DRAM[29351] = 8'b10101;
DRAM[29352] = 8'b110;
DRAM[29353] = 8'b110;
DRAM[29354] = 8'b110;
DRAM[29355] = 8'b110;
DRAM[29356] = 8'b111;
DRAM[29357] = 8'b1000;
DRAM[29358] = 8'b1010;
DRAM[29359] = 8'b1011;
DRAM[29360] = 8'b10101;
DRAM[29361] = 8'b10;
DRAM[29362] = 8'b110;
DRAM[29363] = 8'b10100;
DRAM[29364] = 8'b101000;
DRAM[29365] = 8'b110101;
DRAM[29366] = 8'b1000110;
DRAM[29367] = 8'b1110111;
DRAM[29368] = 8'b10001100;
DRAM[29369] = 8'b10011111;
DRAM[29370] = 8'b10100001;
DRAM[29371] = 8'b10011001;
DRAM[29372] = 8'b10011100;
DRAM[29373] = 8'b10011010;
DRAM[29374] = 8'b10001011;
DRAM[29375] = 8'b10000001;
DRAM[29376] = 8'b10000110;
DRAM[29377] = 8'b10000001;
DRAM[29378] = 8'b1111000;
DRAM[29379] = 8'b1101100;
DRAM[29380] = 8'b1100000;
DRAM[29381] = 8'b1011000;
DRAM[29382] = 8'b1010100;
DRAM[29383] = 8'b1010011;
DRAM[29384] = 8'b1010010;
DRAM[29385] = 8'b1101011;
DRAM[29386] = 8'b1011011;
DRAM[29387] = 8'b1111100;
DRAM[29388] = 8'b10011101;
DRAM[29389] = 8'b10010000;
DRAM[29390] = 8'b10110100;
DRAM[29391] = 8'b11010011;
DRAM[29392] = 8'b11011000;
DRAM[29393] = 8'b11100100;
DRAM[29394] = 8'b11111010;
DRAM[29395] = 8'b11110101;
DRAM[29396] = 8'b11111110;
DRAM[29397] = 8'b11101010;
DRAM[29398] = 8'b11011100;
DRAM[29399] = 8'b11000011;
DRAM[29400] = 8'b10111101;
DRAM[29401] = 8'b10101001;
DRAM[29402] = 8'b10001010;
DRAM[29403] = 8'b10100101;
DRAM[29404] = 8'b10100001;
DRAM[29405] = 8'b10100101;
DRAM[29406] = 8'b10101001;
DRAM[29407] = 8'b10111010;
DRAM[29408] = 8'b10110101;
DRAM[29409] = 8'b10011110;
DRAM[29410] = 8'b10010001;
DRAM[29411] = 8'b1111101;
DRAM[29412] = 8'b1111011;
DRAM[29413] = 8'b10000100;
DRAM[29414] = 8'b1111100;
DRAM[29415] = 8'b10000010;
DRAM[29416] = 8'b1111001;
DRAM[29417] = 8'b1111001;
DRAM[29418] = 8'b1111001;
DRAM[29419] = 8'b1111010;
DRAM[29420] = 8'b1111001;
DRAM[29421] = 8'b1111000;
DRAM[29422] = 8'b1110111;
DRAM[29423] = 8'b1110110;
DRAM[29424] = 8'b1110110;
DRAM[29425] = 8'b1110101;
DRAM[29426] = 8'b1110100;
DRAM[29427] = 8'b1110101;
DRAM[29428] = 8'b1110110;
DRAM[29429] = 8'b1110110;
DRAM[29430] = 8'b1110100;
DRAM[29431] = 8'b1110010;
DRAM[29432] = 8'b1110011;
DRAM[29433] = 8'b1110011;
DRAM[29434] = 8'b1110011;
DRAM[29435] = 8'b1110011;
DRAM[29436] = 8'b1110010;
DRAM[29437] = 8'b1110010;
DRAM[29438] = 8'b1110010;
DRAM[29439] = 8'b1110001;
DRAM[29440] = 8'b10000110;
DRAM[29441] = 8'b10000110;
DRAM[29442] = 8'b10000110;
DRAM[29443] = 8'b10000110;
DRAM[29444] = 8'b10000111;
DRAM[29445] = 8'b10000111;
DRAM[29446] = 8'b10000111;
DRAM[29447] = 8'b10001000;
DRAM[29448] = 8'b10001001;
DRAM[29449] = 8'b10001001;
DRAM[29450] = 8'b10001001;
DRAM[29451] = 8'b10001010;
DRAM[29452] = 8'b10001010;
DRAM[29453] = 8'b10001010;
DRAM[29454] = 8'b10001011;
DRAM[29455] = 8'b10001011;
DRAM[29456] = 8'b10001100;
DRAM[29457] = 8'b10001011;
DRAM[29458] = 8'b10001010;
DRAM[29459] = 8'b10001010;
DRAM[29460] = 8'b10001010;
DRAM[29461] = 8'b10001010;
DRAM[29462] = 8'b10001011;
DRAM[29463] = 8'b10001100;
DRAM[29464] = 8'b10001101;
DRAM[29465] = 8'b10001101;
DRAM[29466] = 8'b10001101;
DRAM[29467] = 8'b10001110;
DRAM[29468] = 8'b10001110;
DRAM[29469] = 8'b10001111;
DRAM[29470] = 8'b10001111;
DRAM[29471] = 8'b10001111;
DRAM[29472] = 8'b10010001;
DRAM[29473] = 8'b10010110;
DRAM[29474] = 8'b10011001;
DRAM[29475] = 8'b10100110;
DRAM[29476] = 8'b10110110;
DRAM[29477] = 8'b10110110;
DRAM[29478] = 8'b10110101;
DRAM[29479] = 8'b11000000;
DRAM[29480] = 8'b10110111;
DRAM[29481] = 8'b10110110;
DRAM[29482] = 8'b10101101;
DRAM[29483] = 8'b10010111;
DRAM[29484] = 8'b10010111;
DRAM[29485] = 8'b10010101;
DRAM[29486] = 8'b10001000;
DRAM[29487] = 8'b10011110;
DRAM[29488] = 8'b10000111;
DRAM[29489] = 8'b10001010;
DRAM[29490] = 8'b10010100;
DRAM[29491] = 8'b10100000;
DRAM[29492] = 8'b10100100;
DRAM[29493] = 8'b10100110;
DRAM[29494] = 8'b10110011;
DRAM[29495] = 8'b11000011;
DRAM[29496] = 8'b10111111;
DRAM[29497] = 8'b11001000;
DRAM[29498] = 8'b11010010;
DRAM[29499] = 8'b11011110;
DRAM[29500] = 8'b11010111;
DRAM[29501] = 8'b11101101;
DRAM[29502] = 8'b11011100;
DRAM[29503] = 8'b11100011;
DRAM[29504] = 8'b11101100;
DRAM[29505] = 8'b11011101;
DRAM[29506] = 8'b11011001;
DRAM[29507] = 8'b11010001;
DRAM[29508] = 8'b10011011;
DRAM[29509] = 8'b11000100;
DRAM[29510] = 8'b10100001;
DRAM[29511] = 8'b10001100;
DRAM[29512] = 8'b1010111;
DRAM[29513] = 8'b1010010;
DRAM[29514] = 8'b1010101;
DRAM[29515] = 8'b1011111;
DRAM[29516] = 8'b1100011;
DRAM[29517] = 8'b1100100;
DRAM[29518] = 8'b1110000;
DRAM[29519] = 8'b10000001;
DRAM[29520] = 8'b10001111;
DRAM[29521] = 8'b10100011;
DRAM[29522] = 8'b10101101;
DRAM[29523] = 8'b10110001;
DRAM[29524] = 8'b10111001;
DRAM[29525] = 8'b10111001;
DRAM[29526] = 8'b10110010;
DRAM[29527] = 8'b10110001;
DRAM[29528] = 8'b10110000;
DRAM[29529] = 8'b10110100;
DRAM[29530] = 8'b11001000;
DRAM[29531] = 8'b11000100;
DRAM[29532] = 8'b10100111;
DRAM[29533] = 8'b10100001;
DRAM[29534] = 8'b10010101;
DRAM[29535] = 8'b1101101;
DRAM[29536] = 8'b1011100;
DRAM[29537] = 8'b10110110;
DRAM[29538] = 8'b11001110;
DRAM[29539] = 8'b11011100;
DRAM[29540] = 8'b10110101;
DRAM[29541] = 8'b1101100;
DRAM[29542] = 8'b1001011;
DRAM[29543] = 8'b100110;
DRAM[29544] = 8'b10010;
DRAM[29545] = 8'b10101;
DRAM[29546] = 8'b1;
DRAM[29547] = 8'b100;
DRAM[29548] = 8'b100101;
DRAM[29549] = 8'b0;
DRAM[29550] = 8'b100000;
DRAM[29551] = 8'b100111;
DRAM[29552] = 8'b0;
DRAM[29553] = 8'b110;
DRAM[29554] = 8'b10;
DRAM[29555] = 8'b10000;
DRAM[29556] = 8'b110011;
DRAM[29557] = 8'b110111;
DRAM[29558] = 8'b110010;
DRAM[29559] = 8'b1000100;
DRAM[29560] = 8'b1000110;
DRAM[29561] = 8'b1001100;
DRAM[29562] = 8'b1011110;
DRAM[29563] = 8'b1110110;
DRAM[29564] = 8'b10000111;
DRAM[29565] = 8'b10001100;
DRAM[29566] = 8'b10010000;
DRAM[29567] = 8'b10010101;
DRAM[29568] = 8'b10011011;
DRAM[29569] = 8'b10100111;
DRAM[29570] = 8'b10100111;
DRAM[29571] = 8'b10100101;
DRAM[29572] = 8'b10101111;
DRAM[29573] = 8'b10110100;
DRAM[29574] = 8'b10110101;
DRAM[29575] = 8'b10111011;
DRAM[29576] = 8'b11001000;
DRAM[29577] = 8'b10111000;
DRAM[29578] = 8'b11000010;
DRAM[29579] = 8'b10111110;
DRAM[29580] = 8'b11000011;
DRAM[29581] = 8'b11001111;
DRAM[29582] = 8'b11001001;
DRAM[29583] = 8'b11000001;
DRAM[29584] = 8'b10111110;
DRAM[29585] = 8'b10111101;
DRAM[29586] = 8'b10111010;
DRAM[29587] = 8'b10110111;
DRAM[29588] = 8'b10110100;
DRAM[29589] = 8'b10110011;
DRAM[29590] = 8'b10110100;
DRAM[29591] = 8'b10110101;
DRAM[29592] = 8'b10100111;
DRAM[29593] = 8'b10101110;
DRAM[29594] = 8'b10101101;
DRAM[29595] = 8'b10100001;
DRAM[29596] = 8'b10110000;
DRAM[29597] = 8'b10010001;
DRAM[29598] = 8'b10011111;
DRAM[29599] = 8'b10110011;
DRAM[29600] = 8'b10101100;
DRAM[29601] = 8'b10000000;
DRAM[29602] = 8'b1101011;
DRAM[29603] = 8'b1000000;
DRAM[29604] = 8'b111011;
DRAM[29605] = 8'b11010;
DRAM[29606] = 8'b10;
DRAM[29607] = 8'b10;
DRAM[29608] = 8'b1001;
DRAM[29609] = 8'b111;
DRAM[29610] = 8'b111;
DRAM[29611] = 8'b1010;
DRAM[29612] = 8'b1011;
DRAM[29613] = 8'b1010;
DRAM[29614] = 8'b1011;
DRAM[29615] = 8'b1101;
DRAM[29616] = 8'b1101;
DRAM[29617] = 8'b1;
DRAM[29618] = 8'b1111;
DRAM[29619] = 8'b100100;
DRAM[29620] = 8'b111101;
DRAM[29621] = 8'b1001001;
DRAM[29622] = 8'b1010011;
DRAM[29623] = 8'b1111100;
DRAM[29624] = 8'b10011110;
DRAM[29625] = 8'b10100111;
DRAM[29626] = 8'b10100000;
DRAM[29627] = 8'b10011000;
DRAM[29628] = 8'b10100001;
DRAM[29629] = 8'b10100110;
DRAM[29630] = 8'b10011100;
DRAM[29631] = 8'b10010110;
DRAM[29632] = 8'b10010100;
DRAM[29633] = 8'b10001110;
DRAM[29634] = 8'b10000011;
DRAM[29635] = 8'b1110011;
DRAM[29636] = 8'b1100011;
DRAM[29637] = 8'b1010111;
DRAM[29638] = 8'b1010010;
DRAM[29639] = 8'b1010000;
DRAM[29640] = 8'b1010001;
DRAM[29641] = 8'b1101100;
DRAM[29642] = 8'b1101010;
DRAM[29643] = 8'b10000100;
DRAM[29644] = 8'b10011000;
DRAM[29645] = 8'b10010111;
DRAM[29646] = 8'b10100010;
DRAM[29647] = 8'b11010100;
DRAM[29648] = 8'b11001100;
DRAM[29649] = 8'b11011010;
DRAM[29650] = 8'b11110101;
DRAM[29651] = 8'b11110110;
DRAM[29652] = 8'b11111111;
DRAM[29653] = 8'b11101110;
DRAM[29654] = 8'b11100010;
DRAM[29655] = 8'b11001100;
DRAM[29656] = 8'b10111111;
DRAM[29657] = 8'b10111010;
DRAM[29658] = 8'b10001111;
DRAM[29659] = 8'b10101001;
DRAM[29660] = 8'b10100101;
DRAM[29661] = 8'b10110000;
DRAM[29662] = 8'b10110101;
DRAM[29663] = 8'b10101111;
DRAM[29664] = 8'b10100010;
DRAM[29665] = 8'b10010001;
DRAM[29666] = 8'b10001101;
DRAM[29667] = 8'b1111111;
DRAM[29668] = 8'b1111110;
DRAM[29669] = 8'b10000100;
DRAM[29670] = 8'b1111001;
DRAM[29671] = 8'b1111011;
DRAM[29672] = 8'b1111010;
DRAM[29673] = 8'b1111010;
DRAM[29674] = 8'b1111010;
DRAM[29675] = 8'b1111001;
DRAM[29676] = 8'b1111001;
DRAM[29677] = 8'b1111000;
DRAM[29678] = 8'b1110111;
DRAM[29679] = 8'b1110111;
DRAM[29680] = 8'b1110111;
DRAM[29681] = 8'b1110110;
DRAM[29682] = 8'b1110101;
DRAM[29683] = 8'b1110110;
DRAM[29684] = 8'b1110111;
DRAM[29685] = 8'b1110111;
DRAM[29686] = 8'b1110101;
DRAM[29687] = 8'b1110011;
DRAM[29688] = 8'b1110100;
DRAM[29689] = 8'b1110100;
DRAM[29690] = 8'b1110011;
DRAM[29691] = 8'b1110011;
DRAM[29692] = 8'b1110011;
DRAM[29693] = 8'b1110010;
DRAM[29694] = 8'b1110010;
DRAM[29695] = 8'b1110010;
DRAM[29696] = 8'b10000110;
DRAM[29697] = 8'b10000111;
DRAM[29698] = 8'b10000111;
DRAM[29699] = 8'b10000111;
DRAM[29700] = 8'b10001000;
DRAM[29701] = 8'b10001000;
DRAM[29702] = 8'b10001000;
DRAM[29703] = 8'b10001000;
DRAM[29704] = 8'b10001001;
DRAM[29705] = 8'b10001001;
DRAM[29706] = 8'b10001010;
DRAM[29707] = 8'b10001010;
DRAM[29708] = 8'b10001010;
DRAM[29709] = 8'b10001011;
DRAM[29710] = 8'b10001011;
DRAM[29711] = 8'b10001011;
DRAM[29712] = 8'b10001100;
DRAM[29713] = 8'b10001100;
DRAM[29714] = 8'b10001011;
DRAM[29715] = 8'b10001010;
DRAM[29716] = 8'b10001010;
DRAM[29717] = 8'b10001011;
DRAM[29718] = 8'b10001100;
DRAM[29719] = 8'b10001100;
DRAM[29720] = 8'b10001101;
DRAM[29721] = 8'b10001101;
DRAM[29722] = 8'b10001110;
DRAM[29723] = 8'b10001110;
DRAM[29724] = 8'b10001110;
DRAM[29725] = 8'b10001110;
DRAM[29726] = 8'b10001111;
DRAM[29727] = 8'b10001111;
DRAM[29728] = 8'b10001110;
DRAM[29729] = 8'b10011011;
DRAM[29730] = 8'b10011011;
DRAM[29731] = 8'b10011000;
DRAM[29732] = 8'b10100011;
DRAM[29733] = 8'b10101100;
DRAM[29734] = 8'b10101110;
DRAM[29735] = 8'b10110010;
DRAM[29736] = 8'b11000000;
DRAM[29737] = 8'b10111110;
DRAM[29738] = 8'b10110010;
DRAM[29739] = 8'b10011011;
DRAM[29740] = 8'b10011100;
DRAM[29741] = 8'b10011001;
DRAM[29742] = 8'b10000110;
DRAM[29743] = 8'b10010100;
DRAM[29744] = 8'b10000111;
DRAM[29745] = 8'b10001010;
DRAM[29746] = 8'b10010110;
DRAM[29747] = 8'b10100100;
DRAM[29748] = 8'b10101000;
DRAM[29749] = 8'b10101001;
DRAM[29750] = 8'b10110110;
DRAM[29751] = 8'b11000101;
DRAM[29752] = 8'b10111100;
DRAM[29753] = 8'b11000011;
DRAM[29754] = 8'b11001100;
DRAM[29755] = 8'b11011010;
DRAM[29756] = 8'b11010110;
DRAM[29757] = 8'b11101110;
DRAM[29758] = 8'b11011011;
DRAM[29759] = 8'b11100001;
DRAM[29760] = 8'b11101001;
DRAM[29761] = 8'b11011010;
DRAM[29762] = 8'b11010100;
DRAM[29763] = 8'b11001011;
DRAM[29764] = 8'b10011100;
DRAM[29765] = 8'b11001000;
DRAM[29766] = 8'b10011111;
DRAM[29767] = 8'b1111111;
DRAM[29768] = 8'b1010111;
DRAM[29769] = 8'b1010111;
DRAM[29770] = 8'b1011010;
DRAM[29771] = 8'b1011111;
DRAM[29772] = 8'b1011111;
DRAM[29773] = 8'b1100010;
DRAM[29774] = 8'b1110000;
DRAM[29775] = 8'b10000000;
DRAM[29776] = 8'b10000010;
DRAM[29777] = 8'b10011000;
DRAM[29778] = 8'b10100101;
DRAM[29779] = 8'b10101001;
DRAM[29780] = 8'b10101101;
DRAM[29781] = 8'b10101010;
DRAM[29782] = 8'b10100111;
DRAM[29783] = 8'b10101110;
DRAM[29784] = 8'b10111100;
DRAM[29785] = 8'b10101101;
DRAM[29786] = 8'b10101110;
DRAM[29787] = 8'b10100111;
DRAM[29788] = 8'b10010110;
DRAM[29789] = 8'b10010110;
DRAM[29790] = 8'b1111111;
DRAM[29791] = 8'b1000110;
DRAM[29792] = 8'b10101110;
DRAM[29793] = 8'b11010111;
DRAM[29794] = 8'b11001110;
DRAM[29795] = 8'b10001011;
DRAM[29796] = 8'b101101;
DRAM[29797] = 8'b101000;
DRAM[29798] = 8'b1010110;
DRAM[29799] = 8'b1001;
DRAM[29800] = 8'b11;
DRAM[29801] = 8'b0;
DRAM[29802] = 8'b1111;
DRAM[29803] = 8'b101100;
DRAM[29804] = 8'b10000000;
DRAM[29805] = 8'b101;
DRAM[29806] = 8'b11001;
DRAM[29807] = 8'b0;
DRAM[29808] = 8'b100;
DRAM[29809] = 8'b11110;
DRAM[29810] = 8'b1110;
DRAM[29811] = 8'b0;
DRAM[29812] = 8'b10111;
DRAM[29813] = 8'b100100;
DRAM[29814] = 8'b100000;
DRAM[29815] = 8'b101101;
DRAM[29816] = 8'b111111;
DRAM[29817] = 8'b1001001;
DRAM[29818] = 8'b1011100;
DRAM[29819] = 8'b1101111;
DRAM[29820] = 8'b1111100;
DRAM[29821] = 8'b10000101;
DRAM[29822] = 8'b10001111;
DRAM[29823] = 8'b10011001;
DRAM[29824] = 8'b10100110;
DRAM[29825] = 8'b10110001;
DRAM[29826] = 8'b10110000;
DRAM[29827] = 8'b10101100;
DRAM[29828] = 8'b10110010;
DRAM[29829] = 8'b10110100;
DRAM[29830] = 8'b10110001;
DRAM[29831] = 8'b10110110;
DRAM[29832] = 8'b11000111;
DRAM[29833] = 8'b10111100;
DRAM[29834] = 8'b11000100;
DRAM[29835] = 8'b11000000;
DRAM[29836] = 8'b10111101;
DRAM[29837] = 8'b11010001;
DRAM[29838] = 8'b11001111;
DRAM[29839] = 8'b11001111;
DRAM[29840] = 8'b11000111;
DRAM[29841] = 8'b11000001;
DRAM[29842] = 8'b10111011;
DRAM[29843] = 8'b10111001;
DRAM[29844] = 8'b10111010;
DRAM[29845] = 8'b10111010;
DRAM[29846] = 8'b10111000;
DRAM[29847] = 8'b10110100;
DRAM[29848] = 8'b10110010;
DRAM[29849] = 8'b11001100;
DRAM[29850] = 8'b10110100;
DRAM[29851] = 8'b10110000;
DRAM[29852] = 8'b11000001;
DRAM[29853] = 8'b10011001;
DRAM[29854] = 8'b10110001;
DRAM[29855] = 8'b10100101;
DRAM[29856] = 8'b10100011;
DRAM[29857] = 8'b10010011;
DRAM[29858] = 8'b1101100;
DRAM[29859] = 8'b1001101;
DRAM[29860] = 8'b1001100;
DRAM[29861] = 8'b11111;
DRAM[29862] = 8'b11101;
DRAM[29863] = 8'b10010;
DRAM[29864] = 8'b1101;
DRAM[29865] = 8'b1000;
DRAM[29866] = 8'b101;
DRAM[29867] = 8'b110;
DRAM[29868] = 8'b100;
DRAM[29869] = 8'b0;
DRAM[29870] = 8'b0;
DRAM[29871] = 8'b1;
DRAM[29872] = 8'b10;
DRAM[29873] = 8'b10100;
DRAM[29874] = 8'b101110;
DRAM[29875] = 8'b110000;
DRAM[29876] = 8'b111000;
DRAM[29877] = 8'b1001010;
DRAM[29878] = 8'b1100011;
DRAM[29879] = 8'b10010010;
DRAM[29880] = 8'b10100100;
DRAM[29881] = 8'b10101101;
DRAM[29882] = 8'b10101000;
DRAM[29883] = 8'b10100000;
DRAM[29884] = 8'b10100101;
DRAM[29885] = 8'b10100110;
DRAM[29886] = 8'b10011101;
DRAM[29887] = 8'b10011010;
DRAM[29888] = 8'b10010011;
DRAM[29889] = 8'b10001011;
DRAM[29890] = 8'b1111110;
DRAM[29891] = 8'b1101111;
DRAM[29892] = 8'b1100000;
DRAM[29893] = 8'b1010101;
DRAM[29894] = 8'b1010000;
DRAM[29895] = 8'b1001110;
DRAM[29896] = 8'b1011010;
DRAM[29897] = 8'b1100110;
DRAM[29898] = 8'b1111101;
DRAM[29899] = 8'b10001110;
DRAM[29900] = 8'b1111111;
DRAM[29901] = 8'b10100000;
DRAM[29902] = 8'b10011001;
DRAM[29903] = 8'b11001100;
DRAM[29904] = 8'b11000100;
DRAM[29905] = 8'b11010000;
DRAM[29906] = 8'b11101110;
DRAM[29907] = 8'b11110010;
DRAM[29908] = 8'b11111111;
DRAM[29909] = 8'b11110000;
DRAM[29910] = 8'b11101000;
DRAM[29911] = 8'b11010110;
DRAM[29912] = 8'b10111010;
DRAM[29913] = 8'b11000011;
DRAM[29914] = 8'b10011101;
DRAM[29915] = 8'b10100110;
DRAM[29916] = 8'b10101000;
DRAM[29917] = 8'b10111001;
DRAM[29918] = 8'b10111101;
DRAM[29919] = 8'b10100011;
DRAM[29920] = 8'b10010100;
DRAM[29921] = 8'b10000111;
DRAM[29922] = 8'b10001000;
DRAM[29923] = 8'b1111111;
DRAM[29924] = 8'b1111111;
DRAM[29925] = 8'b10000100;
DRAM[29926] = 8'b1110111;
DRAM[29927] = 8'b1111001;
DRAM[29928] = 8'b1111100;
DRAM[29929] = 8'b1111011;
DRAM[29930] = 8'b1111010;
DRAM[29931] = 8'b1111001;
DRAM[29932] = 8'b1111000;
DRAM[29933] = 8'b1111000;
DRAM[29934] = 8'b1110111;
DRAM[29935] = 8'b1110111;
DRAM[29936] = 8'b1111000;
DRAM[29937] = 8'b1110111;
DRAM[29938] = 8'b1110110;
DRAM[29939] = 8'b1110111;
DRAM[29940] = 8'b1111000;
DRAM[29941] = 8'b1111000;
DRAM[29942] = 8'b1110101;
DRAM[29943] = 8'b1110011;
DRAM[29944] = 8'b1110100;
DRAM[29945] = 8'b1110100;
DRAM[29946] = 8'b1110100;
DRAM[29947] = 8'b1110011;
DRAM[29948] = 8'b1110011;
DRAM[29949] = 8'b1110011;
DRAM[29950] = 8'b1110010;
DRAM[29951] = 8'b1110010;
DRAM[29952] = 8'b10000111;
DRAM[29953] = 8'b10000111;
DRAM[29954] = 8'b10001000;
DRAM[29955] = 8'b10001000;
DRAM[29956] = 8'b10001000;
DRAM[29957] = 8'b10001001;
DRAM[29958] = 8'b10001001;
DRAM[29959] = 8'b10001001;
DRAM[29960] = 8'b10001010;
DRAM[29961] = 8'b10001010;
DRAM[29962] = 8'b10001010;
DRAM[29963] = 8'b10001010;
DRAM[29964] = 8'b10001011;
DRAM[29965] = 8'b10001011;
DRAM[29966] = 8'b10001011;
DRAM[29967] = 8'b10001100;
DRAM[29968] = 8'b10001100;
DRAM[29969] = 8'b10001100;
DRAM[29970] = 8'b10001011;
DRAM[29971] = 8'b10001011;
DRAM[29972] = 8'b10001011;
DRAM[29973] = 8'b10001011;
DRAM[29974] = 8'b10001100;
DRAM[29975] = 8'b10001100;
DRAM[29976] = 8'b10001110;
DRAM[29977] = 8'b10001110;
DRAM[29978] = 8'b10001110;
DRAM[29979] = 8'b10001110;
DRAM[29980] = 8'b10001110;
DRAM[29981] = 8'b10001110;
DRAM[29982] = 8'b10001110;
DRAM[29983] = 8'b10001110;
DRAM[29984] = 8'b10001001;
DRAM[29985] = 8'b10011001;
DRAM[29986] = 8'b10010111;
DRAM[29987] = 8'b10001111;
DRAM[29988] = 8'b10011001;
DRAM[29989] = 8'b10100101;
DRAM[29990] = 8'b10101000;
DRAM[29991] = 8'b10101001;
DRAM[29992] = 8'b10111011;
DRAM[29993] = 8'b10111001;
DRAM[29994] = 8'b10111000;
DRAM[29995] = 8'b10100100;
DRAM[29996] = 8'b10011110;
DRAM[29997] = 8'b10011011;
DRAM[29998] = 8'b10001001;
DRAM[29999] = 8'b10001110;
DRAM[30000] = 8'b10001010;
DRAM[30001] = 8'b10001101;
DRAM[30002] = 8'b10011000;
DRAM[30003] = 8'b10100101;
DRAM[30004] = 8'b10101000;
DRAM[30005] = 8'b10101000;
DRAM[30006] = 8'b10110100;
DRAM[30007] = 8'b11000011;
DRAM[30008] = 8'b10111001;
DRAM[30009] = 8'b11000000;
DRAM[30010] = 8'b11010000;
DRAM[30011] = 8'b11010110;
DRAM[30012] = 8'b11010111;
DRAM[30013] = 8'b11100111;
DRAM[30014] = 8'b11011100;
DRAM[30015] = 8'b11100000;
DRAM[30016] = 8'b11100111;
DRAM[30017] = 8'b11010011;
DRAM[30018] = 8'b11010111;
DRAM[30019] = 8'b10111111;
DRAM[30020] = 8'b10101101;
DRAM[30021] = 8'b10111001;
DRAM[30022] = 8'b10100110;
DRAM[30023] = 8'b1110010;
DRAM[30024] = 8'b1011111;
DRAM[30025] = 8'b1011101;
DRAM[30026] = 8'b1011001;
DRAM[30027] = 8'b1010110;
DRAM[30028] = 8'b1010111;
DRAM[30029] = 8'b1100000;
DRAM[30030] = 8'b1110000;
DRAM[30031] = 8'b1111110;
DRAM[30032] = 8'b1111000;
DRAM[30033] = 8'b10001100;
DRAM[30034] = 8'b10011000;
DRAM[30035] = 8'b10011100;
DRAM[30036] = 8'b10100000;
DRAM[30037] = 8'b10011101;
DRAM[30038] = 8'b10011111;
DRAM[30039] = 8'b10101011;
DRAM[30040] = 8'b10100101;
DRAM[30041] = 8'b10101111;
DRAM[30042] = 8'b10100000;
DRAM[30043] = 8'b10011001;
DRAM[30044] = 8'b10100011;
DRAM[30045] = 8'b10001110;
DRAM[30046] = 8'b1110100;
DRAM[30047] = 8'b1111100;
DRAM[30048] = 8'b10100001;
DRAM[30049] = 8'b10010111;
DRAM[30050] = 8'b1001010;
DRAM[30051] = 8'b1111;
DRAM[30052] = 8'b10110;
DRAM[30053] = 8'b10010;
DRAM[30054] = 8'b100011;
DRAM[30055] = 8'b10100;
DRAM[30056] = 8'b10001;
DRAM[30057] = 8'b10101;
DRAM[30058] = 8'b0;
DRAM[30059] = 8'b1000;
DRAM[30060] = 8'b11001;
DRAM[30061] = 8'b0;
DRAM[30062] = 8'b10100;
DRAM[30063] = 8'b111;
DRAM[30064] = 8'b1000;
DRAM[30065] = 8'b110001;
DRAM[30066] = 8'b100111;
DRAM[30067] = 8'b110;
DRAM[30068] = 8'b1110;
DRAM[30069] = 8'b10111;
DRAM[30070] = 8'b10010;
DRAM[30071] = 8'b10111;
DRAM[30072] = 8'b111110;
DRAM[30073] = 8'b1001110;
DRAM[30074] = 8'b1100001;
DRAM[30075] = 8'b1101110;
DRAM[30076] = 8'b1111100;
DRAM[30077] = 8'b10001110;
DRAM[30078] = 8'b10011110;
DRAM[30079] = 8'b10100111;
DRAM[30080] = 8'b10101011;
DRAM[30081] = 8'b10110110;
DRAM[30082] = 8'b10110100;
DRAM[30083] = 8'b10101111;
DRAM[30084] = 8'b10110100;
DRAM[30085] = 8'b10110100;
DRAM[30086] = 8'b10110001;
DRAM[30087] = 8'b10110101;
DRAM[30088] = 8'b11000101;
DRAM[30089] = 8'b11000001;
DRAM[30090] = 8'b11000110;
DRAM[30091] = 8'b11000011;
DRAM[30092] = 8'b10111000;
DRAM[30093] = 8'b11010011;
DRAM[30094] = 8'b11010001;
DRAM[30095] = 8'b11010101;
DRAM[30096] = 8'b11001110;
DRAM[30097] = 8'b11001001;
DRAM[30098] = 8'b11000011;
DRAM[30099] = 8'b11000010;
DRAM[30100] = 8'b11000100;
DRAM[30101] = 8'b11000001;
DRAM[30102] = 8'b10111000;
DRAM[30103] = 8'b10110000;
DRAM[30104] = 8'b10111101;
DRAM[30105] = 8'b11011011;
DRAM[30106] = 8'b10110000;
DRAM[30107] = 8'b11000001;
DRAM[30108] = 8'b10110010;
DRAM[30109] = 8'b10101001;
DRAM[30110] = 8'b10101001;
DRAM[30111] = 8'b10010010;
DRAM[30112] = 8'b10001110;
DRAM[30113] = 8'b10011100;
DRAM[30114] = 8'b1110010;
DRAM[30115] = 8'b1011100;
DRAM[30116] = 8'b1011000;
DRAM[30117] = 8'b110011;
DRAM[30118] = 8'b110110;
DRAM[30119] = 8'b101011;
DRAM[30120] = 8'b1111;
DRAM[30121] = 8'b1000;
DRAM[30122] = 8'b110;
DRAM[30123] = 8'b1011;
DRAM[30124] = 8'b1011;
DRAM[30125] = 8'b1000;
DRAM[30126] = 8'b1010;
DRAM[30127] = 8'b10010;
DRAM[30128] = 8'b100100;
DRAM[30129] = 8'b110001;
DRAM[30130] = 8'b111110;
DRAM[30131] = 8'b110101;
DRAM[30132] = 8'b1000100;
DRAM[30133] = 8'b1101000;
DRAM[30134] = 8'b10000001;
DRAM[30135] = 8'b10100100;
DRAM[30136] = 8'b10011011;
DRAM[30137] = 8'b10101000;
DRAM[30138] = 8'b10101000;
DRAM[30139] = 8'b10100001;
DRAM[30140] = 8'b10100000;
DRAM[30141] = 8'b10010111;
DRAM[30142] = 8'b10001010;
DRAM[30143] = 8'b10000111;
DRAM[30144] = 8'b10000110;
DRAM[30145] = 8'b1111101;
DRAM[30146] = 8'b1101111;
DRAM[30147] = 8'b1100010;
DRAM[30148] = 8'b1011010;
DRAM[30149] = 8'b1010110;
DRAM[30150] = 8'b1010011;
DRAM[30151] = 8'b1010010;
DRAM[30152] = 8'b1100101;
DRAM[30153] = 8'b1100101;
DRAM[30154] = 8'b10000011;
DRAM[30155] = 8'b10010001;
DRAM[30156] = 8'b1111101;
DRAM[30157] = 8'b10011001;
DRAM[30158] = 8'b10011001;
DRAM[30159] = 8'b10111011;
DRAM[30160] = 8'b11000001;
DRAM[30161] = 8'b11001001;
DRAM[30162] = 8'b11100011;
DRAM[30163] = 8'b11101011;
DRAM[30164] = 8'b11111111;
DRAM[30165] = 8'b11110010;
DRAM[30166] = 8'b11101110;
DRAM[30167] = 8'b11100000;
DRAM[30168] = 8'b10111001;
DRAM[30169] = 8'b10111110;
DRAM[30170] = 8'b10101110;
DRAM[30171] = 8'b10100011;
DRAM[30172] = 8'b10101101;
DRAM[30173] = 8'b10110111;
DRAM[30174] = 8'b10111000;
DRAM[30175] = 8'b10011100;
DRAM[30176] = 8'b10010000;
DRAM[30177] = 8'b10000011;
DRAM[30178] = 8'b10000011;
DRAM[30179] = 8'b1111001;
DRAM[30180] = 8'b1111001;
DRAM[30181] = 8'b10000001;
DRAM[30182] = 8'b1111001;
DRAM[30183] = 8'b1111110;
DRAM[30184] = 8'b1111101;
DRAM[30185] = 8'b1111100;
DRAM[30186] = 8'b1111011;
DRAM[30187] = 8'b1111001;
DRAM[30188] = 8'b1111000;
DRAM[30189] = 8'b1111000;
DRAM[30190] = 8'b1111000;
DRAM[30191] = 8'b1111000;
DRAM[30192] = 8'b1111001;
DRAM[30193] = 8'b1110111;
DRAM[30194] = 8'b1110111;
DRAM[30195] = 8'b1110111;
DRAM[30196] = 8'b1111001;
DRAM[30197] = 8'b1111000;
DRAM[30198] = 8'b1110110;
DRAM[30199] = 8'b1110100;
DRAM[30200] = 8'b1110101;
DRAM[30201] = 8'b1110100;
DRAM[30202] = 8'b1110100;
DRAM[30203] = 8'b1110100;
DRAM[30204] = 8'b1110011;
DRAM[30205] = 8'b1110011;
DRAM[30206] = 8'b1110011;
DRAM[30207] = 8'b1110011;
DRAM[30208] = 8'b10001000;
DRAM[30209] = 8'b10001000;
DRAM[30210] = 8'b10001000;
DRAM[30211] = 8'b10001001;
DRAM[30212] = 8'b10001001;
DRAM[30213] = 8'b10001001;
DRAM[30214] = 8'b10001010;
DRAM[30215] = 8'b10001010;
DRAM[30216] = 8'b10001010;
DRAM[30217] = 8'b10001010;
DRAM[30218] = 8'b10001010;
DRAM[30219] = 8'b10001011;
DRAM[30220] = 8'b10001011;
DRAM[30221] = 8'b10001011;
DRAM[30222] = 8'b10001100;
DRAM[30223] = 8'b10001100;
DRAM[30224] = 8'b10001101;
DRAM[30225] = 8'b10001100;
DRAM[30226] = 8'b10001100;
DRAM[30227] = 8'b10001011;
DRAM[30228] = 8'b10001011;
DRAM[30229] = 8'b10001100;
DRAM[30230] = 8'b10001100;
DRAM[30231] = 8'b10001101;
DRAM[30232] = 8'b10001110;
DRAM[30233] = 8'b10001110;
DRAM[30234] = 8'b10001110;
DRAM[30235] = 8'b10001110;
DRAM[30236] = 8'b10001110;
DRAM[30237] = 8'b10001110;
DRAM[30238] = 8'b10001110;
DRAM[30239] = 8'b10001110;
DRAM[30240] = 8'b10001100;
DRAM[30241] = 8'b10010101;
DRAM[30242] = 8'b10010100;
DRAM[30243] = 8'b10010011;
DRAM[30244] = 8'b10011100;
DRAM[30245] = 8'b10011111;
DRAM[30246] = 8'b10011110;
DRAM[30247] = 8'b10100011;
DRAM[30248] = 8'b10101110;
DRAM[30249] = 8'b10101111;
DRAM[30250] = 8'b11000000;
DRAM[30251] = 8'b10110011;
DRAM[30252] = 8'b10011111;
DRAM[30253] = 8'b10011110;
DRAM[30254] = 8'b10010101;
DRAM[30255] = 8'b10010011;
DRAM[30256] = 8'b10010000;
DRAM[30257] = 8'b10010010;
DRAM[30258] = 8'b10011100;
DRAM[30259] = 8'b10100111;
DRAM[30260] = 8'b10101000;
DRAM[30261] = 8'b10100111;
DRAM[30262] = 8'b10110010;
DRAM[30263] = 8'b11000001;
DRAM[30264] = 8'b10111000;
DRAM[30265] = 8'b11000001;
DRAM[30266] = 8'b11011100;
DRAM[30267] = 8'b11010101;
DRAM[30268] = 8'b11011000;
DRAM[30269] = 8'b11011011;
DRAM[30270] = 8'b11011011;
DRAM[30271] = 8'b11100010;
DRAM[30272] = 8'b11011101;
DRAM[30273] = 8'b11010011;
DRAM[30274] = 8'b11001110;
DRAM[30275] = 8'b11000010;
DRAM[30276] = 8'b10101101;
DRAM[30277] = 8'b10101001;
DRAM[30278] = 8'b10100001;
DRAM[30279] = 8'b1100111;
DRAM[30280] = 8'b1100000;
DRAM[30281] = 8'b1011110;
DRAM[30282] = 8'b1011010;
DRAM[30283] = 8'b1010111;
DRAM[30284] = 8'b1011011;
DRAM[30285] = 8'b1100101;
DRAM[30286] = 8'b1101111;
DRAM[30287] = 8'b1110101;
DRAM[30288] = 8'b1111010;
DRAM[30289] = 8'b10000111;
DRAM[30290] = 8'b10001110;
DRAM[30291] = 8'b10010010;
DRAM[30292] = 8'b10011001;
DRAM[30293] = 8'b10011010;
DRAM[30294] = 8'b10011110;
DRAM[30295] = 8'b10101100;
DRAM[30296] = 8'b10100011;
DRAM[30297] = 8'b10110110;
DRAM[30298] = 8'b10101110;
DRAM[30299] = 8'b10100101;
DRAM[30300] = 8'b10100111;
DRAM[30301] = 8'b10001101;
DRAM[30302] = 8'b1110011;
DRAM[30303] = 8'b1111100;
DRAM[30304] = 8'b1100011;
DRAM[30305] = 8'b100001;
DRAM[30306] = 8'b111;
DRAM[30307] = 8'b1111;
DRAM[30308] = 8'b100110;
DRAM[30309] = 8'b10011;
DRAM[30310] = 8'b10101;
DRAM[30311] = 8'b1010;
DRAM[30312] = 8'b0;
DRAM[30313] = 8'b100100;
DRAM[30314] = 8'b101;
DRAM[30315] = 8'b11000;
DRAM[30316] = 8'b0;
DRAM[30317] = 8'b10100;
DRAM[30318] = 8'b10101;
DRAM[30319] = 8'b1000;
DRAM[30320] = 8'b110;
DRAM[30321] = 8'b110010;
DRAM[30322] = 8'b110111;
DRAM[30323] = 8'b11011;
DRAM[30324] = 8'b10011;
DRAM[30325] = 8'b10101;
DRAM[30326] = 8'b10101;
DRAM[30327] = 8'b11101;
DRAM[30328] = 8'b110111;
DRAM[30329] = 8'b1001100;
DRAM[30330] = 8'b1011110;
DRAM[30331] = 8'b1101001;
DRAM[30332] = 8'b1111110;
DRAM[30333] = 8'b10011100;
DRAM[30334] = 8'b10101110;
DRAM[30335] = 8'b10101111;
DRAM[30336] = 8'b10101011;
DRAM[30337] = 8'b10110110;
DRAM[30338] = 8'b10110101;
DRAM[30339] = 8'b10110010;
DRAM[30340] = 8'b10111010;
DRAM[30341] = 8'b10111100;
DRAM[30342] = 8'b10111011;
DRAM[30343] = 8'b11000000;
DRAM[30344] = 8'b11001001;
DRAM[30345] = 8'b11001000;
DRAM[30346] = 8'b11001100;
DRAM[30347] = 8'b11001100;
DRAM[30348] = 8'b10111101;
DRAM[30349] = 8'b11011011;
DRAM[30350] = 8'b11010011;
DRAM[30351] = 8'b11010101;
DRAM[30352] = 8'b11011000;
DRAM[30353] = 8'b11010100;
DRAM[30354] = 8'b11001111;
DRAM[30355] = 8'b11001011;
DRAM[30356] = 8'b11001010;
DRAM[30357] = 8'b11001000;
DRAM[30358] = 8'b11000100;
DRAM[30359] = 8'b11000000;
DRAM[30360] = 8'b11001100;
DRAM[30361] = 8'b11000111;
DRAM[30362] = 8'b10111011;
DRAM[30363] = 8'b10111110;
DRAM[30364] = 8'b10101000;
DRAM[30365] = 8'b10110100;
DRAM[30366] = 8'b10011110;
DRAM[30367] = 8'b10010011;
DRAM[30368] = 8'b10101000;
DRAM[30369] = 8'b11000001;
DRAM[30370] = 8'b10011110;
DRAM[30371] = 8'b1110110;
DRAM[30372] = 8'b1011001;
DRAM[30373] = 8'b1000001;
DRAM[30374] = 8'b100101;
DRAM[30375] = 8'b100100;
DRAM[30376] = 8'b101011;
DRAM[30377] = 8'b100011;
DRAM[30378] = 8'b100010;
DRAM[30379] = 8'b101010;
DRAM[30380] = 8'b101110;
DRAM[30381] = 8'b101101;
DRAM[30382] = 8'b110100;
DRAM[30383] = 8'b111110;
DRAM[30384] = 8'b1000001;
DRAM[30385] = 8'b1000000;
DRAM[30386] = 8'b1000101;
DRAM[30387] = 8'b1000111;
DRAM[30388] = 8'b1101010;
DRAM[30389] = 8'b10001111;
DRAM[30390] = 8'b10010100;
DRAM[30391] = 8'b10100001;
DRAM[30392] = 8'b10100000;
DRAM[30393] = 8'b10101100;
DRAM[30394] = 8'b10101011;
DRAM[30395] = 8'b10100101;
DRAM[30396] = 8'b10100101;
DRAM[30397] = 8'b10011110;
DRAM[30398] = 8'b10010100;
DRAM[30399] = 8'b10010100;
DRAM[30400] = 8'b10001101;
DRAM[30401] = 8'b1111111;
DRAM[30402] = 8'b1101110;
DRAM[30403] = 8'b1100011;
DRAM[30404] = 8'b1011111;
DRAM[30405] = 8'b1011111;
DRAM[30406] = 8'b1011100;
DRAM[30407] = 8'b1011010;
DRAM[30408] = 8'b1100101;
DRAM[30409] = 8'b1101100;
DRAM[30410] = 8'b10000000;
DRAM[30411] = 8'b10011001;
DRAM[30412] = 8'b10101100;
DRAM[30413] = 8'b10000111;
DRAM[30414] = 8'b10011010;
DRAM[30415] = 8'b10011111;
DRAM[30416] = 8'b11000001;
DRAM[30417] = 8'b11000100;
DRAM[30418] = 8'b11011010;
DRAM[30419] = 8'b11100010;
DRAM[30420] = 8'b11111011;
DRAM[30421] = 8'b11110010;
DRAM[30422] = 8'b11110010;
DRAM[30423] = 8'b11100111;
DRAM[30424] = 8'b11000011;
DRAM[30425] = 8'b10110101;
DRAM[30426] = 8'b10111111;
DRAM[30427] = 8'b10100100;
DRAM[30428] = 8'b10110101;
DRAM[30429] = 8'b10101001;
DRAM[30430] = 8'b10100100;
DRAM[30431] = 8'b10010110;
DRAM[30432] = 8'b10001100;
DRAM[30433] = 8'b10000000;
DRAM[30434] = 8'b10000010;
DRAM[30435] = 8'b1111000;
DRAM[30436] = 8'b1111001;
DRAM[30437] = 8'b10000001;
DRAM[30438] = 8'b1111010;
DRAM[30439] = 8'b10000000;
DRAM[30440] = 8'b1111111;
DRAM[30441] = 8'b1111101;
DRAM[30442] = 8'b1111011;
DRAM[30443] = 8'b1111001;
DRAM[30444] = 8'b1111000;
DRAM[30445] = 8'b1110111;
DRAM[30446] = 8'b1111000;
DRAM[30447] = 8'b1111000;
DRAM[30448] = 8'b1111001;
DRAM[30449] = 8'b1111000;
DRAM[30450] = 8'b1110111;
DRAM[30451] = 8'b1111000;
DRAM[30452] = 8'b1111001;
DRAM[30453] = 8'b1111001;
DRAM[30454] = 8'b1110111;
DRAM[30455] = 8'b1110101;
DRAM[30456] = 8'b1110101;
DRAM[30457] = 8'b1110101;
DRAM[30458] = 8'b1110100;
DRAM[30459] = 8'b1110100;
DRAM[30460] = 8'b1110100;
DRAM[30461] = 8'b1110011;
DRAM[30462] = 8'b1110011;
DRAM[30463] = 8'b1110011;
DRAM[30464] = 8'b10001000;
DRAM[30465] = 8'b10001000;
DRAM[30466] = 8'b10001001;
DRAM[30467] = 8'b10001001;
DRAM[30468] = 8'b10001001;
DRAM[30469] = 8'b10001010;
DRAM[30470] = 8'b10001010;
DRAM[30471] = 8'b10001010;
DRAM[30472] = 8'b10001010;
DRAM[30473] = 8'b10001010;
DRAM[30474] = 8'b10001010;
DRAM[30475] = 8'b10001011;
DRAM[30476] = 8'b10001011;
DRAM[30477] = 8'b10001100;
DRAM[30478] = 8'b10001100;
DRAM[30479] = 8'b10001100;
DRAM[30480] = 8'b10001101;
DRAM[30481] = 8'b10001100;
DRAM[30482] = 8'b10001100;
DRAM[30483] = 8'b10001011;
DRAM[30484] = 8'b10001011;
DRAM[30485] = 8'b10001100;
DRAM[30486] = 8'b10001100;
DRAM[30487] = 8'b10001101;
DRAM[30488] = 8'b10001110;
DRAM[30489] = 8'b10001110;
DRAM[30490] = 8'b10001110;
DRAM[30491] = 8'b10001110;
DRAM[30492] = 8'b10001110;
DRAM[30493] = 8'b10001110;
DRAM[30494] = 8'b10001110;
DRAM[30495] = 8'b10001110;
DRAM[30496] = 8'b10010011;
DRAM[30497] = 8'b10010011;
DRAM[30498] = 8'b10010010;
DRAM[30499] = 8'b10011011;
DRAM[30500] = 8'b10100100;
DRAM[30501] = 8'b10011010;
DRAM[30502] = 8'b10010100;
DRAM[30503] = 8'b10011111;
DRAM[30504] = 8'b10101000;
DRAM[30505] = 8'b10101101;
DRAM[30506] = 8'b11001101;
DRAM[30507] = 8'b11000011;
DRAM[30508] = 8'b10100110;
DRAM[30509] = 8'b10100110;
DRAM[30510] = 8'b10100100;
DRAM[30511] = 8'b10100001;
DRAM[30512] = 8'b10010110;
DRAM[30513] = 8'b10011000;
DRAM[30514] = 8'b10100000;
DRAM[30515] = 8'b10101001;
DRAM[30516] = 8'b10101010;
DRAM[30517] = 8'b10101000;
DRAM[30518] = 8'b10110010;
DRAM[30519] = 8'b11000000;
DRAM[30520] = 8'b10110111;
DRAM[30521] = 8'b11000011;
DRAM[30522] = 8'b11101000;
DRAM[30523] = 8'b11010110;
DRAM[30524] = 8'b11011000;
DRAM[30525] = 8'b11010001;
DRAM[30526] = 8'b11011010;
DRAM[30527] = 8'b11100100;
DRAM[30528] = 8'b11010001;
DRAM[30529] = 8'b11011001;
DRAM[30530] = 8'b10111100;
DRAM[30531] = 8'b11010001;
DRAM[30532] = 8'b10011011;
DRAM[30533] = 8'b10100100;
DRAM[30534] = 8'b10010011;
DRAM[30535] = 8'b1100001;
DRAM[30536] = 8'b1011010;
DRAM[30537] = 8'b1011101;
DRAM[30538] = 8'b1011111;
DRAM[30539] = 8'b1100001;
DRAM[30540] = 8'b1100111;
DRAM[30541] = 8'b1101110;
DRAM[30542] = 8'b1101110;
DRAM[30543] = 8'b1101010;
DRAM[30544] = 8'b1111110;
DRAM[30545] = 8'b10000101;
DRAM[30546] = 8'b10000101;
DRAM[30547] = 8'b10001010;
DRAM[30548] = 8'b10010110;
DRAM[30549] = 8'b10011010;
DRAM[30550] = 8'b10011101;
DRAM[30551] = 8'b10101001;
DRAM[30552] = 8'b10100100;
DRAM[30553] = 8'b10011001;
DRAM[30554] = 8'b10100000;
DRAM[30555] = 8'b10100101;
DRAM[30556] = 8'b10100100;
DRAM[30557] = 8'b10101110;
DRAM[30558] = 8'b10010000;
DRAM[30559] = 8'b1001010;
DRAM[30560] = 8'b110001;
DRAM[30561] = 8'b101001;
DRAM[30562] = 8'b11101;
DRAM[30563] = 8'b0;
DRAM[30564] = 8'b11001;
DRAM[30565] = 8'b10001;
DRAM[30566] = 8'b1001;
DRAM[30567] = 8'b10011;
DRAM[30568] = 8'b10111;
DRAM[30569] = 8'b0;
DRAM[30570] = 8'b11;
DRAM[30571] = 8'b10001;
DRAM[30572] = 8'b100111;
DRAM[30573] = 8'b0;
DRAM[30574] = 8'b10001;
DRAM[30575] = 8'b0;
DRAM[30576] = 8'b11;
DRAM[30577] = 8'b101010;
DRAM[30578] = 8'b111001;
DRAM[30579] = 8'b101000;
DRAM[30580] = 8'b11001;
DRAM[30581] = 8'b10110;
DRAM[30582] = 8'b100000;
DRAM[30583] = 8'b110001;
DRAM[30584] = 8'b101000;
DRAM[30585] = 8'b111111;
DRAM[30586] = 8'b1010000;
DRAM[30587] = 8'b1011100;
DRAM[30588] = 8'b1111000;
DRAM[30589] = 8'b10011111;
DRAM[30590] = 8'b10110000;
DRAM[30591] = 8'b10101010;
DRAM[30592] = 8'b10101010;
DRAM[30593] = 8'b10110110;
DRAM[30594] = 8'b10110111;
DRAM[30595] = 8'b10110110;
DRAM[30596] = 8'b11000000;
DRAM[30597] = 8'b11000110;
DRAM[30598] = 8'b11000111;
DRAM[30599] = 8'b11001101;
DRAM[30600] = 8'b11001111;
DRAM[30601] = 8'b11001111;
DRAM[30602] = 8'b11010010;
DRAM[30603] = 8'b11010101;
DRAM[30604] = 8'b11000101;
DRAM[30605] = 8'b11100011;
DRAM[30606] = 8'b11010101;
DRAM[30607] = 8'b11010010;
DRAM[30608] = 8'b11100001;
DRAM[30609] = 8'b11011101;
DRAM[30610] = 8'b11010110;
DRAM[30611] = 8'b11001110;
DRAM[30612] = 8'b11001011;
DRAM[30613] = 8'b11001110;
DRAM[30614] = 8'b11010101;
DRAM[30615] = 8'b11011011;
DRAM[30616] = 8'b11011110;
DRAM[30617] = 8'b10101101;
DRAM[30618] = 8'b11010011;
DRAM[30619] = 8'b10110010;
DRAM[30620] = 8'b10110010;
DRAM[30621] = 8'b10111001;
DRAM[30622] = 8'b10100100;
DRAM[30623] = 8'b10100110;
DRAM[30624] = 8'b10101110;
DRAM[30625] = 8'b11001011;
DRAM[30626] = 8'b10111100;
DRAM[30627] = 8'b10001000;
DRAM[30628] = 8'b1100011;
DRAM[30629] = 8'b1100000;
DRAM[30630] = 8'b101101;
DRAM[30631] = 8'b111100;
DRAM[30632] = 8'b111111;
DRAM[30633] = 8'b110101;
DRAM[30634] = 8'b110001;
DRAM[30635] = 8'b110101;
DRAM[30636] = 8'b110110;
DRAM[30637] = 8'b110011;
DRAM[30638] = 8'b111000;
DRAM[30639] = 8'b1000011;
DRAM[30640] = 8'b110011;
DRAM[30641] = 8'b111101;
DRAM[30642] = 8'b1010101;
DRAM[30643] = 8'b1100101;
DRAM[30644] = 8'b10000010;
DRAM[30645] = 8'b10010101;
DRAM[30646] = 8'b10001110;
DRAM[30647] = 8'b10011001;
DRAM[30648] = 8'b10100000;
DRAM[30649] = 8'b10100101;
DRAM[30650] = 8'b10011111;
DRAM[30651] = 8'b10011010;
DRAM[30652] = 8'b10100001;
DRAM[30653] = 8'b10100011;
DRAM[30654] = 8'b10100010;
DRAM[30655] = 8'b10101001;
DRAM[30656] = 8'b10100001;
DRAM[30657] = 8'b10010000;
DRAM[30658] = 8'b1111010;
DRAM[30659] = 8'b1101101;
DRAM[30660] = 8'b1101001;
DRAM[30661] = 8'b1101000;
DRAM[30662] = 8'b1100100;
DRAM[30663] = 8'b1011111;
DRAM[30664] = 8'b1011110;
DRAM[30665] = 8'b1110100;
DRAM[30666] = 8'b1111101;
DRAM[30667] = 8'b10100100;
DRAM[30668] = 8'b11100100;
DRAM[30669] = 8'b1111010;
DRAM[30670] = 8'b10011011;
DRAM[30671] = 8'b10000111;
DRAM[30672] = 8'b11000011;
DRAM[30673] = 8'b11000001;
DRAM[30674] = 8'b11010100;
DRAM[30675] = 8'b11011101;
DRAM[30676] = 8'b11111000;
DRAM[30677] = 8'b11110010;
DRAM[30678] = 8'b11110101;
DRAM[30679] = 8'b11101011;
DRAM[30680] = 8'b11010001;
DRAM[30681] = 8'b10101111;
DRAM[30682] = 8'b11001010;
DRAM[30683] = 8'b10101001;
DRAM[30684] = 8'b10111011;
DRAM[30685] = 8'b10011001;
DRAM[30686] = 8'b10010000;
DRAM[30687] = 8'b10001111;
DRAM[30688] = 8'b10000101;
DRAM[30689] = 8'b1111101;
DRAM[30690] = 8'b10000011;
DRAM[30691] = 8'b1111101;
DRAM[30692] = 8'b1111110;
DRAM[30693] = 8'b10000011;
DRAM[30694] = 8'b1111000;
DRAM[30695] = 8'b1111100;
DRAM[30696] = 8'b1111111;
DRAM[30697] = 8'b1111110;
DRAM[30698] = 8'b1111011;
DRAM[30699] = 8'b1111001;
DRAM[30700] = 8'b1111000;
DRAM[30701] = 8'b1110111;
DRAM[30702] = 8'b1111000;
DRAM[30703] = 8'b1111000;
DRAM[30704] = 8'b1111001;
DRAM[30705] = 8'b1111000;
DRAM[30706] = 8'b1111000;
DRAM[30707] = 8'b1111000;
DRAM[30708] = 8'b1111001;
DRAM[30709] = 8'b1111001;
DRAM[30710] = 8'b1110111;
DRAM[30711] = 8'b1110101;
DRAM[30712] = 8'b1110101;
DRAM[30713] = 8'b1110101;
DRAM[30714] = 8'b1110101;
DRAM[30715] = 8'b1110100;
DRAM[30716] = 8'b1110100;
DRAM[30717] = 8'b1110011;
DRAM[30718] = 8'b1110011;
DRAM[30719] = 8'b1110011;
DRAM[30720] = 8'b10001001;
DRAM[30721] = 8'b10001001;
DRAM[30722] = 8'b10001001;
DRAM[30723] = 8'b10001001;
DRAM[30724] = 8'b10001001;
DRAM[30725] = 8'b10001001;
DRAM[30726] = 8'b10001001;
DRAM[30727] = 8'b10001001;
DRAM[30728] = 8'b10001001;
DRAM[30729] = 8'b10001010;
DRAM[30730] = 8'b10001011;
DRAM[30731] = 8'b10001100;
DRAM[30732] = 8'b10001100;
DRAM[30733] = 8'b10001100;
DRAM[30734] = 8'b10001011;
DRAM[30735] = 8'b10001011;
DRAM[30736] = 8'b10001110;
DRAM[30737] = 8'b10001101;
DRAM[30738] = 8'b10001101;
DRAM[30739] = 8'b10001101;
DRAM[30740] = 8'b10001101;
DRAM[30741] = 8'b10001110;
DRAM[30742] = 8'b10001111;
DRAM[30743] = 8'b10010000;
DRAM[30744] = 8'b10010000;
DRAM[30745] = 8'b10010000;
DRAM[30746] = 8'b10010000;
DRAM[30747] = 8'b10010001;
DRAM[30748] = 8'b10010001;
DRAM[30749] = 8'b10010010;
DRAM[30750] = 8'b10010010;
DRAM[30751] = 8'b10010010;
DRAM[30752] = 8'b10010001;
DRAM[30753] = 8'b10010010;
DRAM[30754] = 8'b10010011;
DRAM[30755] = 8'b10010101;
DRAM[30756] = 8'b10010111;
DRAM[30757] = 8'b10011001;
DRAM[30758] = 8'b10011011;
DRAM[30759] = 8'b10011011;
DRAM[30760] = 8'b10011100;
DRAM[30761] = 8'b10111011;
DRAM[30762] = 8'b10110101;
DRAM[30763] = 8'b10111011;
DRAM[30764] = 8'b10111100;
DRAM[30765] = 8'b10101110;
DRAM[30766] = 8'b10110001;
DRAM[30767] = 8'b10100001;
DRAM[30768] = 8'b10100110;
DRAM[30769] = 8'b10100110;
DRAM[30770] = 8'b10100110;
DRAM[30771] = 8'b10011011;
DRAM[30772] = 8'b10100100;
DRAM[30773] = 8'b10010111;
DRAM[30774] = 8'b10111110;
DRAM[30775] = 8'b11001001;
DRAM[30776] = 8'b11001000;
DRAM[30777] = 8'b11100000;
DRAM[30778] = 8'b11100010;
DRAM[30779] = 8'b11010110;
DRAM[30780] = 8'b11011101;
DRAM[30781] = 8'b11001110;
DRAM[30782] = 8'b11101011;
DRAM[30783] = 8'b11010110;
DRAM[30784] = 8'b11011100;
DRAM[30785] = 8'b11001101;
DRAM[30786] = 8'b10111011;
DRAM[30787] = 8'b10111011;
DRAM[30788] = 8'b10011010;
DRAM[30789] = 8'b10100000;
DRAM[30790] = 8'b10000011;
DRAM[30791] = 8'b1100010;
DRAM[30792] = 8'b1011000;
DRAM[30793] = 8'b1010110;
DRAM[30794] = 8'b1011001;
DRAM[30795] = 8'b1100001;
DRAM[30796] = 8'b1101010;
DRAM[30797] = 8'b1110001;
DRAM[30798] = 8'b1111010;
DRAM[30799] = 8'b10000010;
DRAM[30800] = 8'b10010001;
DRAM[30801] = 8'b10010110;
DRAM[30802] = 8'b10011000;
DRAM[30803] = 8'b10010001;
DRAM[30804] = 8'b10000111;
DRAM[30805] = 8'b10000111;
DRAM[30806] = 8'b10010010;
DRAM[30807] = 8'b10011110;
DRAM[30808] = 8'b10100110;
DRAM[30809] = 8'b10100011;
DRAM[30810] = 8'b10100100;
DRAM[30811] = 8'b10100010;
DRAM[30812] = 8'b10100010;
DRAM[30813] = 8'b10100011;
DRAM[30814] = 8'b10001011;
DRAM[30815] = 8'b1100010;
DRAM[30816] = 8'b1001001;
DRAM[30817] = 8'b101000;
DRAM[30818] = 8'b101100;
DRAM[30819] = 8'b10001;
DRAM[30820] = 8'b10010;
DRAM[30821] = 8'b100011;
DRAM[30822] = 8'b101;
DRAM[30823] = 8'b1110;
DRAM[30824] = 8'b101;
DRAM[30825] = 8'b1000;
DRAM[30826] = 8'b1010;
DRAM[30827] = 8'b1010;
DRAM[30828] = 8'b1100;
DRAM[30829] = 8'b1101;
DRAM[30830] = 8'b1000;
DRAM[30831] = 8'b0;
DRAM[30832] = 8'b0;
DRAM[30833] = 8'b111100;
DRAM[30834] = 8'b111111;
DRAM[30835] = 8'b100011;
DRAM[30836] = 8'b11000;
DRAM[30837] = 8'b11101;
DRAM[30838] = 8'b110100;
DRAM[30839] = 8'b111111;
DRAM[30840] = 8'b111111;
DRAM[30841] = 8'b1011101;
DRAM[30842] = 8'b1100100;
DRAM[30843] = 8'b1110000;
DRAM[30844] = 8'b10010100;
DRAM[30845] = 8'b10100000;
DRAM[30846] = 8'b10100010;
DRAM[30847] = 8'b10111001;
DRAM[30848] = 8'b10110010;
DRAM[30849] = 8'b10101110;
DRAM[30850] = 8'b10110011;
DRAM[30851] = 8'b10111111;
DRAM[30852] = 8'b11001000;
DRAM[30853] = 8'b11000111;
DRAM[30854] = 8'b11000110;
DRAM[30855] = 8'b11000111;
DRAM[30856] = 8'b11010010;
DRAM[30857] = 8'b11011011;
DRAM[30858] = 8'b11011001;
DRAM[30859] = 8'b11010011;
DRAM[30860] = 8'b11010100;
DRAM[30861] = 8'b11010010;
DRAM[30862] = 8'b11010110;
DRAM[30863] = 8'b11100100;
DRAM[30864] = 8'b11101011;
DRAM[30865] = 8'b11011010;
DRAM[30866] = 8'b11001111;
DRAM[30867] = 8'b11010010;
DRAM[30868] = 8'b11010110;
DRAM[30869] = 8'b11010110;
DRAM[30870] = 8'b11011010;
DRAM[30871] = 8'b11100011;
DRAM[30872] = 8'b11001010;
DRAM[30873] = 8'b11001011;
DRAM[30874] = 8'b11010011;
DRAM[30875] = 8'b10111101;
DRAM[30876] = 8'b10111110;
DRAM[30877] = 8'b10101011;
DRAM[30878] = 8'b10110000;
DRAM[30879] = 8'b10101000;
DRAM[30880] = 8'b10100111;
DRAM[30881] = 8'b11001010;
DRAM[30882] = 8'b11001001;
DRAM[30883] = 8'b10011111;
DRAM[30884] = 8'b1110000;
DRAM[30885] = 8'b1000110;
DRAM[30886] = 8'b110111;
DRAM[30887] = 8'b1001000;
DRAM[30888] = 8'b1100001;
DRAM[30889] = 8'b1010010;
DRAM[30890] = 8'b111101;
DRAM[30891] = 8'b111101;
DRAM[30892] = 8'b111110;
DRAM[30893] = 8'b1100001;
DRAM[30894] = 8'b1001010;
DRAM[30895] = 8'b1000100;
DRAM[30896] = 8'b1011101;
DRAM[30897] = 8'b1010111;
DRAM[30898] = 8'b1100110;
DRAM[30899] = 8'b10001001;
DRAM[30900] = 8'b10011100;
DRAM[30901] = 8'b10011010;
DRAM[30902] = 8'b10011100;
DRAM[30903] = 8'b10100111;
DRAM[30904] = 8'b10011001;
DRAM[30905] = 8'b10011111;
DRAM[30906] = 8'b10100101;
DRAM[30907] = 8'b10101010;
DRAM[30908] = 8'b10101101;
DRAM[30909] = 8'b10101011;
DRAM[30910] = 8'b10011110;
DRAM[30911] = 8'b10010000;
DRAM[30912] = 8'b10001000;
DRAM[30913] = 8'b10000011;
DRAM[30914] = 8'b10000110;
DRAM[30915] = 8'b10000000;
DRAM[30916] = 8'b1101000;
DRAM[30917] = 8'b1011011;
DRAM[30918] = 8'b1011100;
DRAM[30919] = 8'b1011100;
DRAM[30920] = 8'b1101101;
DRAM[30921] = 8'b1111111;
DRAM[30922] = 8'b1111101;
DRAM[30923] = 8'b10011111;
DRAM[30924] = 8'b11010100;
DRAM[30925] = 8'b10111000;
DRAM[30926] = 8'b10000110;
DRAM[30927] = 8'b10010001;
DRAM[30928] = 8'b10100011;
DRAM[30929] = 8'b10110000;
DRAM[30930] = 8'b10111011;
DRAM[30931] = 8'b11110111;
DRAM[30932] = 8'b11110000;
DRAM[30933] = 8'b11110100;
DRAM[30934] = 8'b11110111;
DRAM[30935] = 8'b11100110;
DRAM[30936] = 8'b11011111;
DRAM[30937] = 8'b10111011;
DRAM[30938] = 8'b11000101;
DRAM[30939] = 8'b10111010;
DRAM[30940] = 8'b10100100;
DRAM[30941] = 8'b10100000;
DRAM[30942] = 8'b10001101;
DRAM[30943] = 8'b10001000;
DRAM[30944] = 8'b10000000;
DRAM[30945] = 8'b10000000;
DRAM[30946] = 8'b10000000;
DRAM[30947] = 8'b1111111;
DRAM[30948] = 8'b1111111;
DRAM[30949] = 8'b1111110;
DRAM[30950] = 8'b1111110;
DRAM[30951] = 8'b1111110;
DRAM[30952] = 8'b1111011;
DRAM[30953] = 8'b1111100;
DRAM[30954] = 8'b1111100;
DRAM[30955] = 8'b1111100;
DRAM[30956] = 8'b1111100;
DRAM[30957] = 8'b1111011;
DRAM[30958] = 8'b1111010;
DRAM[30959] = 8'b1111001;
DRAM[30960] = 8'b1111001;
DRAM[30961] = 8'b1111001;
DRAM[30962] = 8'b1111000;
DRAM[30963] = 8'b1111000;
DRAM[30964] = 8'b1111000;
DRAM[30965] = 8'b1110111;
DRAM[30966] = 8'b1110111;
DRAM[30967] = 8'b1110111;
DRAM[30968] = 8'b1110110;
DRAM[30969] = 8'b1110110;
DRAM[30970] = 8'b1110101;
DRAM[30971] = 8'b1110100;
DRAM[30972] = 8'b1110100;
DRAM[30973] = 8'b1110011;
DRAM[30974] = 8'b1110010;
DRAM[30975] = 8'b1110010;
DRAM[30976] = 8'b10001001;
DRAM[30977] = 8'b10001001;
DRAM[30978] = 8'b10001001;
DRAM[30979] = 8'b10001001;
DRAM[30980] = 8'b10001001;
DRAM[30981] = 8'b10001001;
DRAM[30982] = 8'b10001001;
DRAM[30983] = 8'b10001001;
DRAM[30984] = 8'b10001001;
DRAM[30985] = 8'b10001010;
DRAM[30986] = 8'b10001011;
DRAM[30987] = 8'b10001100;
DRAM[30988] = 8'b10001100;
DRAM[30989] = 8'b10001100;
DRAM[30990] = 8'b10001100;
DRAM[30991] = 8'b10001011;
DRAM[30992] = 8'b10001110;
DRAM[30993] = 8'b10001110;
DRAM[30994] = 8'b10001101;
DRAM[30995] = 8'b10001101;
DRAM[30996] = 8'b10001110;
DRAM[30997] = 8'b10001110;
DRAM[30998] = 8'b10001111;
DRAM[30999] = 8'b10010000;
DRAM[31000] = 8'b10001111;
DRAM[31001] = 8'b10001111;
DRAM[31002] = 8'b10001111;
DRAM[31003] = 8'b10010000;
DRAM[31004] = 8'b10010000;
DRAM[31005] = 8'b10010000;
DRAM[31006] = 8'b10010001;
DRAM[31007] = 8'b10010001;
DRAM[31008] = 8'b10010001;
DRAM[31009] = 8'b10010010;
DRAM[31010] = 8'b10010011;
DRAM[31011] = 8'b10010100;
DRAM[31012] = 8'b10010110;
DRAM[31013] = 8'b10010111;
DRAM[31014] = 8'b10011000;
DRAM[31015] = 8'b10011001;
DRAM[31016] = 8'b10010111;
DRAM[31017] = 8'b10101001;
DRAM[31018] = 8'b10101010;
DRAM[31019] = 8'b10111000;
DRAM[31020] = 8'b10111001;
DRAM[31021] = 8'b10110000;
DRAM[31022] = 8'b10110110;
DRAM[31023] = 8'b10100101;
DRAM[31024] = 8'b10101011;
DRAM[31025] = 8'b10101000;
DRAM[31026] = 8'b10100101;
DRAM[31027] = 8'b10100000;
DRAM[31028] = 8'b10101101;
DRAM[31029] = 8'b10100011;
DRAM[31030] = 8'b11000011;
DRAM[31031] = 8'b11000111;
DRAM[31032] = 8'b11000111;
DRAM[31033] = 8'b11001111;
DRAM[31034] = 8'b11100001;
DRAM[31035] = 8'b11001100;
DRAM[31036] = 8'b11010111;
DRAM[31037] = 8'b11011011;
DRAM[31038] = 8'b11100101;
DRAM[31039] = 8'b11011110;
DRAM[31040] = 8'b11010010;
DRAM[31041] = 8'b11000111;
DRAM[31042] = 8'b10111000;
DRAM[31043] = 8'b10111000;
DRAM[31044] = 8'b10011011;
DRAM[31045] = 8'b10011110;
DRAM[31046] = 8'b10000010;
DRAM[31047] = 8'b1100010;
DRAM[31048] = 8'b1100100;
DRAM[31049] = 8'b1011111;
DRAM[31050] = 8'b1011101;
DRAM[31051] = 8'b1100001;
DRAM[31052] = 8'b1100101;
DRAM[31053] = 8'b1101010;
DRAM[31054] = 8'b1110010;
DRAM[31055] = 8'b1111010;
DRAM[31056] = 8'b1111011;
DRAM[31057] = 8'b10000011;
DRAM[31058] = 8'b10001110;
DRAM[31059] = 8'b10010101;
DRAM[31060] = 8'b10010110;
DRAM[31061] = 8'b10010011;
DRAM[31062] = 8'b10010001;
DRAM[31063] = 8'b10010000;
DRAM[31064] = 8'b10101010;
DRAM[31065] = 8'b10101010;
DRAM[31066] = 8'b10110000;
DRAM[31067] = 8'b10110010;
DRAM[31068] = 8'b10110011;
DRAM[31069] = 8'b10111000;
DRAM[31070] = 8'b10100110;
DRAM[31071] = 8'b10000010;
DRAM[31072] = 8'b1010011;
DRAM[31073] = 8'b1000001;
DRAM[31074] = 8'b110110;
DRAM[31075] = 8'b100100;
DRAM[31076] = 8'b1111;
DRAM[31077] = 8'b100;
DRAM[31078] = 8'b1000;
DRAM[31079] = 8'b100000;
DRAM[31080] = 8'b1000;
DRAM[31081] = 8'b1010;
DRAM[31082] = 8'b111;
DRAM[31083] = 8'b10;
DRAM[31084] = 8'b0;
DRAM[31085] = 8'b11;
DRAM[31086] = 8'b100;
DRAM[31087] = 8'b11;
DRAM[31088] = 8'b1000;
DRAM[31089] = 8'b111100;
DRAM[31090] = 8'b110001;
DRAM[31091] = 8'b10111;
DRAM[31092] = 8'b10101;
DRAM[31093] = 8'b10110;
DRAM[31094] = 8'b101110;
DRAM[31095] = 8'b1000111;
DRAM[31096] = 8'b1001010;
DRAM[31097] = 8'b1011010;
DRAM[31098] = 8'b1101000;
DRAM[31099] = 8'b10001000;
DRAM[31100] = 8'b10110011;
DRAM[31101] = 8'b10111010;
DRAM[31102] = 8'b10101001;
DRAM[31103] = 8'b10100101;
DRAM[31104] = 8'b10110111;
DRAM[31105] = 8'b10110101;
DRAM[31106] = 8'b10111000;
DRAM[31107] = 8'b11000000;
DRAM[31108] = 8'b11000101;
DRAM[31109] = 8'b11001010;
DRAM[31110] = 8'b11010100;
DRAM[31111] = 8'b11011110;
DRAM[31112] = 8'b11011000;
DRAM[31113] = 8'b11011110;
DRAM[31114] = 8'b11011001;
DRAM[31115] = 8'b11010111;
DRAM[31116] = 8'b11011101;
DRAM[31117] = 8'b11011101;
DRAM[31118] = 8'b11011010;
DRAM[31119] = 8'b11100001;
DRAM[31120] = 8'b11101110;
DRAM[31121] = 8'b11100001;
DRAM[31122] = 8'b11011010;
DRAM[31123] = 8'b11011111;
DRAM[31124] = 8'b11100011;
DRAM[31125] = 8'b11100001;
DRAM[31126] = 8'b11100011;
DRAM[31127] = 8'b11101001;
DRAM[31128] = 8'b11010111;
DRAM[31129] = 8'b11010100;
DRAM[31130] = 8'b11001111;
DRAM[31131] = 8'b11001111;
DRAM[31132] = 8'b11000010;
DRAM[31133] = 8'b10110111;
DRAM[31134] = 8'b10110011;
DRAM[31135] = 8'b10111011;
DRAM[31136] = 8'b10111011;
DRAM[31137] = 8'b11001011;
DRAM[31138] = 8'b11001001;
DRAM[31139] = 8'b10110011;
DRAM[31140] = 8'b10010111;
DRAM[31141] = 8'b1110110;
DRAM[31142] = 8'b1011011;
DRAM[31143] = 8'b1010001;
DRAM[31144] = 8'b1001110;
DRAM[31145] = 8'b1100110;
DRAM[31146] = 8'b1110010;
DRAM[31147] = 8'b1011111;
DRAM[31148] = 8'b110110;
DRAM[31149] = 8'b1000101;
DRAM[31150] = 8'b1001101;
DRAM[31151] = 8'b1101111;
DRAM[31152] = 8'b1101000;
DRAM[31153] = 8'b1110010;
DRAM[31154] = 8'b1111001;
DRAM[31155] = 8'b1111100;
DRAM[31156] = 8'b10001001;
DRAM[31157] = 8'b10011110;
DRAM[31158] = 8'b10101011;
DRAM[31159] = 8'b10101101;
DRAM[31160] = 8'b10100110;
DRAM[31161] = 8'b10100101;
DRAM[31162] = 8'b10100000;
DRAM[31163] = 8'b10011101;
DRAM[31164] = 8'b10011111;
DRAM[31165] = 8'b10100010;
DRAM[31166] = 8'b10011110;
DRAM[31167] = 8'b10011000;
DRAM[31168] = 8'b10001111;
DRAM[31169] = 8'b10001001;
DRAM[31170] = 8'b10001011;
DRAM[31171] = 8'b10000100;
DRAM[31172] = 8'b1101110;
DRAM[31173] = 8'b1100100;
DRAM[31174] = 8'b1101000;
DRAM[31175] = 8'b1101001;
DRAM[31176] = 8'b1100011;
DRAM[31177] = 8'b1111001;
DRAM[31178] = 8'b1111111;
DRAM[31179] = 8'b10011101;
DRAM[31180] = 8'b11010000;
DRAM[31181] = 8'b11000011;
DRAM[31182] = 8'b10001111;
DRAM[31183] = 8'b1111110;
DRAM[31184] = 8'b10100000;
DRAM[31185] = 8'b10110000;
DRAM[31186] = 8'b10110100;
DRAM[31187] = 8'b11100101;
DRAM[31188] = 8'b11101011;
DRAM[31189] = 8'b11110101;
DRAM[31190] = 8'b11110111;
DRAM[31191] = 8'b11101010;
DRAM[31192] = 8'b11100100;
DRAM[31193] = 8'b11000010;
DRAM[31194] = 8'b11000011;
DRAM[31195] = 8'b10110100;
DRAM[31196] = 8'b10011101;
DRAM[31197] = 8'b10011000;
DRAM[31198] = 8'b10001001;
DRAM[31199] = 8'b10000100;
DRAM[31200] = 8'b10000000;
DRAM[31201] = 8'b10000000;
DRAM[31202] = 8'b10000000;
DRAM[31203] = 8'b1111111;
DRAM[31204] = 8'b1111111;
DRAM[31205] = 8'b1111111;
DRAM[31206] = 8'b1111110;
DRAM[31207] = 8'b1111110;
DRAM[31208] = 8'b1111101;
DRAM[31209] = 8'b1111101;
DRAM[31210] = 8'b1111101;
DRAM[31211] = 8'b1111101;
DRAM[31212] = 8'b1111101;
DRAM[31213] = 8'b1111100;
DRAM[31214] = 8'b1111011;
DRAM[31215] = 8'b1111011;
DRAM[31216] = 8'b1111001;
DRAM[31217] = 8'b1111000;
DRAM[31218] = 8'b1111000;
DRAM[31219] = 8'b1111000;
DRAM[31220] = 8'b1110111;
DRAM[31221] = 8'b1110111;
DRAM[31222] = 8'b1110111;
DRAM[31223] = 8'b1110110;
DRAM[31224] = 8'b1110111;
DRAM[31225] = 8'b1110111;
DRAM[31226] = 8'b1110111;
DRAM[31227] = 8'b1110110;
DRAM[31228] = 8'b1110101;
DRAM[31229] = 8'b1110100;
DRAM[31230] = 8'b1110100;
DRAM[31231] = 8'b1110011;
DRAM[31232] = 8'b10001010;
DRAM[31233] = 8'b10001010;
DRAM[31234] = 8'b10001010;
DRAM[31235] = 8'b10001010;
DRAM[31236] = 8'b10001010;
DRAM[31237] = 8'b10001010;
DRAM[31238] = 8'b10001010;
DRAM[31239] = 8'b10001010;
DRAM[31240] = 8'b10001010;
DRAM[31241] = 8'b10001011;
DRAM[31242] = 8'b10001100;
DRAM[31243] = 8'b10001100;
DRAM[31244] = 8'b10001101;
DRAM[31245] = 8'b10001101;
DRAM[31246] = 8'b10001100;
DRAM[31247] = 8'b10001100;
DRAM[31248] = 8'b10001110;
DRAM[31249] = 8'b10001110;
DRAM[31250] = 8'b10001101;
DRAM[31251] = 8'b10001101;
DRAM[31252] = 8'b10001110;
DRAM[31253] = 8'b10001111;
DRAM[31254] = 8'b10010000;
DRAM[31255] = 8'b10010000;
DRAM[31256] = 8'b10001110;
DRAM[31257] = 8'b10001110;
DRAM[31258] = 8'b10001111;
DRAM[31259] = 8'b10001111;
DRAM[31260] = 8'b10001111;
DRAM[31261] = 8'b10010000;
DRAM[31262] = 8'b10010000;
DRAM[31263] = 8'b10010000;
DRAM[31264] = 8'b10010001;
DRAM[31265] = 8'b10010010;
DRAM[31266] = 8'b10010010;
DRAM[31267] = 8'b10010011;
DRAM[31268] = 8'b10010100;
DRAM[31269] = 8'b10010101;
DRAM[31270] = 8'b10010101;
DRAM[31271] = 8'b10010110;
DRAM[31272] = 8'b10011100;
DRAM[31273] = 8'b10011100;
DRAM[31274] = 8'b10100110;
DRAM[31275] = 8'b10111011;
DRAM[31276] = 8'b10110110;
DRAM[31277] = 8'b10110010;
DRAM[31278] = 8'b10111111;
DRAM[31279] = 8'b10110001;
DRAM[31280] = 8'b10101111;
DRAM[31281] = 8'b10101001;
DRAM[31282] = 8'b10011111;
DRAM[31283] = 8'b10100000;
DRAM[31284] = 8'b10101110;
DRAM[31285] = 8'b10101000;
DRAM[31286] = 8'b10111110;
DRAM[31287] = 8'b10111101;
DRAM[31288] = 8'b11001010;
DRAM[31289] = 8'b11000100;
DRAM[31290] = 8'b11011111;
DRAM[31291] = 8'b11000110;
DRAM[31292] = 8'b11010010;
DRAM[31293] = 8'b11100100;
DRAM[31294] = 8'b11011011;
DRAM[31295] = 8'b11011111;
DRAM[31296] = 8'b11000101;
DRAM[31297] = 8'b10111110;
DRAM[31298] = 8'b10110011;
DRAM[31299] = 8'b10110001;
DRAM[31300] = 8'b10011100;
DRAM[31301] = 8'b10011010;
DRAM[31302] = 8'b10000000;
DRAM[31303] = 8'b1100010;
DRAM[31304] = 8'b1101101;
DRAM[31305] = 8'b1100110;
DRAM[31306] = 8'b1100001;
DRAM[31307] = 8'b1100010;
DRAM[31308] = 8'b1100100;
DRAM[31309] = 8'b1100111;
DRAM[31310] = 8'b1101110;
DRAM[31311] = 8'b1110110;
DRAM[31312] = 8'b1111001;
DRAM[31313] = 8'b1111010;
DRAM[31314] = 8'b10000000;
DRAM[31315] = 8'b10001011;
DRAM[31316] = 8'b10010110;
DRAM[31317] = 8'b10011101;
DRAM[31318] = 8'b10011101;
DRAM[31319] = 8'b10011010;
DRAM[31320] = 8'b10011011;
DRAM[31321] = 8'b10011111;
DRAM[31322] = 8'b10101010;
DRAM[31323] = 8'b10101111;
DRAM[31324] = 8'b10110001;
DRAM[31325] = 8'b10111010;
DRAM[31326] = 8'b10110010;
DRAM[31327] = 8'b10011000;
DRAM[31328] = 8'b1111001;
DRAM[31329] = 8'b1011000;
DRAM[31330] = 8'b101101;
DRAM[31331] = 8'b101010;
DRAM[31332] = 8'b11111;
DRAM[31333] = 8'b100;
DRAM[31334] = 8'b111;
DRAM[31335] = 8'b1000;
DRAM[31336] = 8'b100;
DRAM[31337] = 8'b1001;
DRAM[31338] = 8'b1100;
DRAM[31339] = 8'b1001;
DRAM[31340] = 8'b111;
DRAM[31341] = 8'b111;
DRAM[31342] = 8'b101;
DRAM[31343] = 8'b1;
DRAM[31344] = 8'b1111;
DRAM[31345] = 8'b110100;
DRAM[31346] = 8'b11111;
DRAM[31347] = 8'b10101;
DRAM[31348] = 8'b100010;
DRAM[31349] = 8'b11010;
DRAM[31350] = 8'b101110;
DRAM[31351] = 8'b1010111;
DRAM[31352] = 8'b1011010;
DRAM[31353] = 8'b1100111;
DRAM[31354] = 8'b10000001;
DRAM[31355] = 8'b10011111;
DRAM[31356] = 8'b10110000;
DRAM[31357] = 8'b10101111;
DRAM[31358] = 8'b10101100;
DRAM[31359] = 8'b10101111;
DRAM[31360] = 8'b10111101;
DRAM[31361] = 8'b11000000;
DRAM[31362] = 8'b11000111;
DRAM[31363] = 8'b11001100;
DRAM[31364] = 8'b11001111;
DRAM[31365] = 8'b11010100;
DRAM[31366] = 8'b11100010;
DRAM[31367] = 8'b11101111;
DRAM[31368] = 8'b11100001;
DRAM[31369] = 8'b11100010;
DRAM[31370] = 8'b11011011;
DRAM[31371] = 8'b11011100;
DRAM[31372] = 8'b11101000;
DRAM[31373] = 8'b11101000;
DRAM[31374] = 8'b11100000;
DRAM[31375] = 8'b11100000;
DRAM[31376] = 8'b11101100;
DRAM[31377] = 8'b11100011;
DRAM[31378] = 8'b11100000;
DRAM[31379] = 8'b11100111;
DRAM[31380] = 8'b11101011;
DRAM[31381] = 8'b11101000;
DRAM[31382] = 8'b11100111;
DRAM[31383] = 8'b11101011;
DRAM[31384] = 8'b11100111;
DRAM[31385] = 8'b11100001;
DRAM[31386] = 8'b11010010;
DRAM[31387] = 8'b11100100;
DRAM[31388] = 8'b11001101;
DRAM[31389] = 8'b11001010;
DRAM[31390] = 8'b11000000;
DRAM[31391] = 8'b11010011;
DRAM[31392] = 8'b11000110;
DRAM[31393] = 8'b11000110;
DRAM[31394] = 8'b11001011;
DRAM[31395] = 8'b11000111;
DRAM[31396] = 8'b10110110;
DRAM[31397] = 8'b10100011;
DRAM[31398] = 8'b10001100;
DRAM[31399] = 8'b1110011;
DRAM[31400] = 8'b1011010;
DRAM[31401] = 8'b1100010;
DRAM[31402] = 8'b1101110;
DRAM[31403] = 8'b1110010;
DRAM[31404] = 8'b1101100;
DRAM[31405] = 8'b1110110;
DRAM[31406] = 8'b1011000;
DRAM[31407] = 8'b1001110;
DRAM[31408] = 8'b1110101;
DRAM[31409] = 8'b10000111;
DRAM[31410] = 8'b10010000;
DRAM[31411] = 8'b10001010;
DRAM[31412] = 8'b10001011;
DRAM[31413] = 8'b10011000;
DRAM[31414] = 8'b10011100;
DRAM[31415] = 8'b10010101;
DRAM[31416] = 8'b10100000;
DRAM[31417] = 8'b10100100;
DRAM[31418] = 8'b10100111;
DRAM[31419] = 8'b10101001;
DRAM[31420] = 8'b10101100;
DRAM[31421] = 8'b10101101;
DRAM[31422] = 8'b10100110;
DRAM[31423] = 8'b10011101;
DRAM[31424] = 8'b10010000;
DRAM[31425] = 8'b10000111;
DRAM[31426] = 8'b10000111;
DRAM[31427] = 8'b10000000;
DRAM[31428] = 8'b1101100;
DRAM[31429] = 8'b1100101;
DRAM[31430] = 8'b1101100;
DRAM[31431] = 8'b1101111;
DRAM[31432] = 8'b1110011;
DRAM[31433] = 8'b10001001;
DRAM[31434] = 8'b10011000;
DRAM[31435] = 8'b10110010;
DRAM[31436] = 8'b11011011;
DRAM[31437] = 8'b11011100;
DRAM[31438] = 8'b10100111;
DRAM[31439] = 8'b1110110;
DRAM[31440] = 8'b10011000;
DRAM[31441] = 8'b10101110;
DRAM[31442] = 8'b10101101;
DRAM[31443] = 8'b11001101;
DRAM[31444] = 8'b11100010;
DRAM[31445] = 8'b11110010;
DRAM[31446] = 8'b11110010;
DRAM[31447] = 8'b11101101;
DRAM[31448] = 8'b11101101;
DRAM[31449] = 8'b11001111;
DRAM[31450] = 8'b11000011;
DRAM[31451] = 8'b10101011;
DRAM[31452] = 8'b10010100;
DRAM[31453] = 8'b10010000;
DRAM[31454] = 8'b10000110;
DRAM[31455] = 8'b10000011;
DRAM[31456] = 8'b10000000;
DRAM[31457] = 8'b10000000;
DRAM[31458] = 8'b10000000;
DRAM[31459] = 8'b10000000;
DRAM[31460] = 8'b1111111;
DRAM[31461] = 8'b1111111;
DRAM[31462] = 8'b1111111;
DRAM[31463] = 8'b1111110;
DRAM[31464] = 8'b1111110;
DRAM[31465] = 8'b1111110;
DRAM[31466] = 8'b1111110;
DRAM[31467] = 8'b1111110;
DRAM[31468] = 8'b1111101;
DRAM[31469] = 8'b1111101;
DRAM[31470] = 8'b1111100;
DRAM[31471] = 8'b1111100;
DRAM[31472] = 8'b1111001;
DRAM[31473] = 8'b1111001;
DRAM[31474] = 8'b1111001;
DRAM[31475] = 8'b1111000;
DRAM[31476] = 8'b1111000;
DRAM[31477] = 8'b1111000;
DRAM[31478] = 8'b1110111;
DRAM[31479] = 8'b1110111;
DRAM[31480] = 8'b1111001;
DRAM[31481] = 8'b1111000;
DRAM[31482] = 8'b1111000;
DRAM[31483] = 8'b1110111;
DRAM[31484] = 8'b1110110;
DRAM[31485] = 8'b1110101;
DRAM[31486] = 8'b1110101;
DRAM[31487] = 8'b1110101;
DRAM[31488] = 8'b10001011;
DRAM[31489] = 8'b10001011;
DRAM[31490] = 8'b10001011;
DRAM[31491] = 8'b10001011;
DRAM[31492] = 8'b10001011;
DRAM[31493] = 8'b10001011;
DRAM[31494] = 8'b10001011;
DRAM[31495] = 8'b10001011;
DRAM[31496] = 8'b10001011;
DRAM[31497] = 8'b10001011;
DRAM[31498] = 8'b10001100;
DRAM[31499] = 8'b10001101;
DRAM[31500] = 8'b10001110;
DRAM[31501] = 8'b10001110;
DRAM[31502] = 8'b10001101;
DRAM[31503] = 8'b10001101;
DRAM[31504] = 8'b10001111;
DRAM[31505] = 8'b10001110;
DRAM[31506] = 8'b10001110;
DRAM[31507] = 8'b10001110;
DRAM[31508] = 8'b10001110;
DRAM[31509] = 8'b10001111;
DRAM[31510] = 8'b10010000;
DRAM[31511] = 8'b10010001;
DRAM[31512] = 8'b10001111;
DRAM[31513] = 8'b10001111;
DRAM[31514] = 8'b10010000;
DRAM[31515] = 8'b10010000;
DRAM[31516] = 8'b10010000;
DRAM[31517] = 8'b10010001;
DRAM[31518] = 8'b10010001;
DRAM[31519] = 8'b10010001;
DRAM[31520] = 8'b10010010;
DRAM[31521] = 8'b10010010;
DRAM[31522] = 8'b10010010;
DRAM[31523] = 8'b10010010;
DRAM[31524] = 8'b10010011;
DRAM[31525] = 8'b10010011;
DRAM[31526] = 8'b10010011;
DRAM[31527] = 8'b10010011;
DRAM[31528] = 8'b10100010;
DRAM[31529] = 8'b10010100;
DRAM[31530] = 8'b10100110;
DRAM[31531] = 8'b10111001;
DRAM[31532] = 8'b10101011;
DRAM[31533] = 8'b10101100;
DRAM[31534] = 8'b11000010;
DRAM[31535] = 8'b10111100;
DRAM[31536] = 8'b10110011;
DRAM[31537] = 8'b10101101;
DRAM[31538] = 8'b10011110;
DRAM[31539] = 8'b10100010;
DRAM[31540] = 8'b10101001;
DRAM[31541] = 8'b10100110;
DRAM[31542] = 8'b10111000;
DRAM[31543] = 8'b10111001;
DRAM[31544] = 8'b11001101;
DRAM[31545] = 8'b11001011;
DRAM[31546] = 8'b11011000;
DRAM[31547] = 8'b11001011;
DRAM[31548] = 8'b11010100;
DRAM[31549] = 8'b11100001;
DRAM[31550] = 8'b11010101;
DRAM[31551] = 8'b11010000;
DRAM[31552] = 8'b10111100;
DRAM[31553] = 8'b10111001;
DRAM[31554] = 8'b10101111;
DRAM[31555] = 8'b10100101;
DRAM[31556] = 8'b10011000;
DRAM[31557] = 8'b10010011;
DRAM[31558] = 8'b1111101;
DRAM[31559] = 8'b1100101;
DRAM[31560] = 8'b1101100;
DRAM[31561] = 8'b1100111;
DRAM[31562] = 8'b1100100;
DRAM[31563] = 8'b1100110;
DRAM[31564] = 8'b1101001;
DRAM[31565] = 8'b1101100;
DRAM[31566] = 8'b1110011;
DRAM[31567] = 8'b1111010;
DRAM[31568] = 8'b1111111;
DRAM[31569] = 8'b1111110;
DRAM[31570] = 8'b10000001;
DRAM[31571] = 8'b10001011;
DRAM[31572] = 8'b10011010;
DRAM[31573] = 8'b10100101;
DRAM[31574] = 8'b10101000;
DRAM[31575] = 8'b10101000;
DRAM[31576] = 8'b10100101;
DRAM[31577] = 8'b10101001;
DRAM[31578] = 8'b10110001;
DRAM[31579] = 8'b10110010;
DRAM[31580] = 8'b10101111;
DRAM[31581] = 8'b10110111;
DRAM[31582] = 8'b10110110;
DRAM[31583] = 8'b10100110;
DRAM[31584] = 8'b10011001;
DRAM[31585] = 8'b1101010;
DRAM[31586] = 8'b111101;
DRAM[31587] = 8'b110101;
DRAM[31588] = 8'b111000;
DRAM[31589] = 8'b101010;
DRAM[31590] = 8'b10100;
DRAM[31591] = 8'b11;
DRAM[31592] = 8'b0;
DRAM[31593] = 8'b0;
DRAM[31594] = 8'b0;
DRAM[31595] = 8'b0;
DRAM[31596] = 8'b0;
DRAM[31597] = 8'b11;
DRAM[31598] = 8'b1;
DRAM[31599] = 8'b0;
DRAM[31600] = 8'b10;
DRAM[31601] = 8'b11111;
DRAM[31602] = 8'b1110;
DRAM[31603] = 8'b11001;
DRAM[31604] = 8'b110100;
DRAM[31605] = 8'b100100;
DRAM[31606] = 8'b110001;
DRAM[31607] = 8'b1100001;
DRAM[31608] = 8'b1101110;
DRAM[31609] = 8'b1111011;
DRAM[31610] = 8'b10011100;
DRAM[31611] = 8'b10110011;
DRAM[31612] = 8'b10101011;
DRAM[31613] = 8'b10100010;
DRAM[31614] = 8'b10101011;
DRAM[31615] = 8'b10110110;
DRAM[31616] = 8'b11000001;
DRAM[31617] = 8'b11001010;
DRAM[31618] = 8'b11010111;
DRAM[31619] = 8'b11011111;
DRAM[31620] = 8'b11100010;
DRAM[31621] = 8'b11100011;
DRAM[31622] = 8'b11100111;
DRAM[31623] = 8'b11101101;
DRAM[31624] = 8'b11101000;
DRAM[31625] = 8'b11101000;
DRAM[31626] = 8'b11100001;
DRAM[31627] = 8'b11100001;
DRAM[31628] = 8'b11101101;
DRAM[31629] = 8'b11101101;
DRAM[31630] = 8'b11100110;
DRAM[31631] = 8'b11100110;
DRAM[31632] = 8'b11101011;
DRAM[31633] = 8'b11100101;
DRAM[31634] = 8'b11100101;
DRAM[31635] = 8'b11101011;
DRAM[31636] = 8'b11101110;
DRAM[31637] = 8'b11101100;
DRAM[31638] = 8'b11101100;
DRAM[31639] = 8'b11101110;
DRAM[31640] = 8'b11110000;
DRAM[31641] = 8'b11101101;
DRAM[31642] = 8'b11100100;
DRAM[31643] = 8'b11101101;
DRAM[31644] = 8'b11011110;
DRAM[31645] = 8'b11011100;
DRAM[31646] = 8'b11010110;
DRAM[31647] = 8'b11100001;
DRAM[31648] = 8'b11010000;
DRAM[31649] = 8'b11001011;
DRAM[31650] = 8'b11010101;
DRAM[31651] = 8'b11010100;
DRAM[31652] = 8'b10111011;
DRAM[31653] = 8'b10101111;
DRAM[31654] = 8'b10100111;
DRAM[31655] = 8'b10010100;
DRAM[31656] = 8'b1111001;
DRAM[31657] = 8'b1110010;
DRAM[31658] = 8'b1110010;
DRAM[31659] = 8'b1101010;
DRAM[31660] = 8'b1101111;
DRAM[31661] = 8'b10000000;
DRAM[31662] = 8'b1110000;
DRAM[31663] = 8'b1101010;
DRAM[31664] = 8'b1110100;
DRAM[31665] = 8'b1111010;
DRAM[31666] = 8'b10001001;
DRAM[31667] = 8'b10011001;
DRAM[31668] = 8'b10011110;
DRAM[31669] = 8'b10011011;
DRAM[31670] = 8'b10011011;
DRAM[31671] = 8'b10011111;
DRAM[31672] = 8'b10010011;
DRAM[31673] = 8'b10011011;
DRAM[31674] = 8'b10100011;
DRAM[31675] = 8'b10101000;
DRAM[31676] = 8'b10101010;
DRAM[31677] = 8'b10100111;
DRAM[31678] = 8'b10011011;
DRAM[31679] = 8'b10010000;
DRAM[31680] = 8'b10010001;
DRAM[31681] = 8'b10000110;
DRAM[31682] = 8'b10000011;
DRAM[31683] = 8'b1111011;
DRAM[31684] = 8'b1101001;
DRAM[31685] = 8'b1100011;
DRAM[31686] = 8'b1101100;
DRAM[31687] = 8'b1110000;
DRAM[31688] = 8'b1110101;
DRAM[31689] = 8'b10000100;
DRAM[31690] = 8'b10011110;
DRAM[31691] = 8'b10111110;
DRAM[31692] = 8'b11011100;
DRAM[31693] = 8'b11100010;
DRAM[31694] = 8'b10111000;
DRAM[31695] = 8'b1111111;
DRAM[31696] = 8'b10001001;
DRAM[31697] = 8'b10100110;
DRAM[31698] = 8'b10101011;
DRAM[31699] = 8'b10111011;
DRAM[31700] = 8'b11011001;
DRAM[31701] = 8'b11101010;
DRAM[31702] = 8'b11101010;
DRAM[31703] = 8'b11101110;
DRAM[31704] = 8'b11110011;
DRAM[31705] = 8'b11011100;
DRAM[31706] = 8'b11000010;
DRAM[31707] = 8'b10100011;
DRAM[31708] = 8'b10001110;
DRAM[31709] = 8'b10001001;
DRAM[31710] = 8'b10000110;
DRAM[31711] = 8'b10000101;
DRAM[31712] = 8'b10000001;
DRAM[31713] = 8'b10000001;
DRAM[31714] = 8'b10000000;
DRAM[31715] = 8'b10000000;
DRAM[31716] = 8'b10000000;
DRAM[31717] = 8'b1111111;
DRAM[31718] = 8'b1111111;
DRAM[31719] = 8'b1111111;
DRAM[31720] = 8'b1111110;
DRAM[31721] = 8'b1111110;
DRAM[31722] = 8'b1111101;
DRAM[31723] = 8'b1111100;
DRAM[31724] = 8'b1111100;
DRAM[31725] = 8'b1111100;
DRAM[31726] = 8'b1111100;
DRAM[31727] = 8'b1111100;
DRAM[31728] = 8'b1111011;
DRAM[31729] = 8'b1111011;
DRAM[31730] = 8'b1111011;
DRAM[31731] = 8'b1111010;
DRAM[31732] = 8'b1111010;
DRAM[31733] = 8'b1111001;
DRAM[31734] = 8'b1111001;
DRAM[31735] = 8'b1111001;
DRAM[31736] = 8'b1111001;
DRAM[31737] = 8'b1111000;
DRAM[31738] = 8'b1111000;
DRAM[31739] = 8'b1110111;
DRAM[31740] = 8'b1110110;
DRAM[31741] = 8'b1110101;
DRAM[31742] = 8'b1110101;
DRAM[31743] = 8'b1110100;
DRAM[31744] = 8'b10001011;
DRAM[31745] = 8'b10001011;
DRAM[31746] = 8'b10001011;
DRAM[31747] = 8'b10001011;
DRAM[31748] = 8'b10001011;
DRAM[31749] = 8'b10001011;
DRAM[31750] = 8'b10001011;
DRAM[31751] = 8'b10001011;
DRAM[31752] = 8'b10001100;
DRAM[31753] = 8'b10001100;
DRAM[31754] = 8'b10001101;
DRAM[31755] = 8'b10001110;
DRAM[31756] = 8'b10001110;
DRAM[31757] = 8'b10001110;
DRAM[31758] = 8'b10001110;
DRAM[31759] = 8'b10001110;
DRAM[31760] = 8'b10001111;
DRAM[31761] = 8'b10001111;
DRAM[31762] = 8'b10001110;
DRAM[31763] = 8'b10001110;
DRAM[31764] = 8'b10001111;
DRAM[31765] = 8'b10001111;
DRAM[31766] = 8'b10010000;
DRAM[31767] = 8'b10010001;
DRAM[31768] = 8'b10010001;
DRAM[31769] = 8'b10010001;
DRAM[31770] = 8'b10010001;
DRAM[31771] = 8'b10010010;
DRAM[31772] = 8'b10010010;
DRAM[31773] = 8'b10010010;
DRAM[31774] = 8'b10010011;
DRAM[31775] = 8'b10010011;
DRAM[31776] = 8'b10010011;
DRAM[31777] = 8'b10010011;
DRAM[31778] = 8'b10010011;
DRAM[31779] = 8'b10010011;
DRAM[31780] = 8'b10010011;
DRAM[31781] = 8'b10010011;
DRAM[31782] = 8'b10010011;
DRAM[31783] = 8'b10010011;
DRAM[31784] = 8'b10011110;
DRAM[31785] = 8'b10001101;
DRAM[31786] = 8'b10100010;
DRAM[31787] = 8'b10101101;
DRAM[31788] = 8'b10011011;
DRAM[31789] = 8'b10100011;
DRAM[31790] = 8'b10111101;
DRAM[31791] = 8'b11000011;
DRAM[31792] = 8'b10110101;
DRAM[31793] = 8'b10110100;
DRAM[31794] = 8'b10100010;
DRAM[31795] = 8'b10101000;
DRAM[31796] = 8'b10100101;
DRAM[31797] = 8'b10100111;
DRAM[31798] = 8'b10111011;
DRAM[31799] = 8'b11000100;
DRAM[31800] = 8'b11001011;
DRAM[31801] = 8'b11011000;
DRAM[31802] = 8'b11001101;
DRAM[31803] = 8'b11010111;
DRAM[31804] = 8'b11011001;
DRAM[31805] = 8'b11010111;
DRAM[31806] = 8'b11010101;
DRAM[31807] = 8'b10111111;
DRAM[31808] = 8'b10111000;
DRAM[31809] = 8'b10110110;
DRAM[31810] = 8'b10101011;
DRAM[31811] = 8'b10011000;
DRAM[31812] = 8'b10010101;
DRAM[31813] = 8'b10001011;
DRAM[31814] = 8'b1111011;
DRAM[31815] = 8'b1101010;
DRAM[31816] = 8'b1101010;
DRAM[31817] = 8'b1100111;
DRAM[31818] = 8'b1101000;
DRAM[31819] = 8'b1101101;
DRAM[31820] = 8'b1110001;
DRAM[31821] = 8'b1110011;
DRAM[31822] = 8'b1111000;
DRAM[31823] = 8'b1111110;
DRAM[31824] = 8'b1111100;
DRAM[31825] = 8'b10000010;
DRAM[31826] = 8'b10001101;
DRAM[31827] = 8'b10011010;
DRAM[31828] = 8'b10100100;
DRAM[31829] = 8'b10101001;
DRAM[31830] = 8'b10101000;
DRAM[31831] = 8'b10100110;
DRAM[31832] = 8'b10101111;
DRAM[31833] = 8'b10101111;
DRAM[31834] = 8'b10110011;
DRAM[31835] = 8'b10101111;
DRAM[31836] = 8'b10100110;
DRAM[31837] = 8'b10101101;
DRAM[31838] = 8'b10110010;
DRAM[31839] = 8'b10101001;
DRAM[31840] = 8'b10011110;
DRAM[31841] = 8'b10000001;
DRAM[31842] = 8'b1111000;
DRAM[31843] = 8'b1001111;
DRAM[31844] = 8'b111101;
DRAM[31845] = 8'b1000010;
DRAM[31846] = 8'b100111;
DRAM[31847] = 8'b101100;
DRAM[31848] = 8'b11010;
DRAM[31849] = 8'b10010;
DRAM[31850] = 8'b111;
DRAM[31851] = 8'b1;
DRAM[31852] = 8'b1000;
DRAM[31853] = 8'b10001;
DRAM[31854] = 8'b10010;
DRAM[31855] = 8'b1100;
DRAM[31856] = 8'b0;
DRAM[31857] = 8'b10011;
DRAM[31858] = 8'b1000;
DRAM[31859] = 8'b11101;
DRAM[31860] = 8'b111001;
DRAM[31861] = 8'b101011;
DRAM[31862] = 8'b111011;
DRAM[31863] = 8'b1101000;
DRAM[31864] = 8'b1111110;
DRAM[31865] = 8'b10001010;
DRAM[31866] = 8'b10101010;
DRAM[31867] = 8'b11000001;
DRAM[31868] = 8'b10111100;
DRAM[31869] = 8'b10110000;
DRAM[31870] = 8'b10101110;
DRAM[31871] = 8'b10101101;
DRAM[31872] = 8'b11000101;
DRAM[31873] = 8'b11001110;
DRAM[31874] = 8'b11011011;
DRAM[31875] = 8'b11100101;
DRAM[31876] = 8'b11101010;
DRAM[31877] = 8'b11101100;
DRAM[31878] = 8'b11101100;
DRAM[31879] = 8'b11101010;
DRAM[31880] = 8'b11101100;
DRAM[31881] = 8'b11101111;
DRAM[31882] = 8'b11101000;
DRAM[31883] = 8'b11100101;
DRAM[31884] = 8'b11101100;
DRAM[31885] = 8'b11101100;
DRAM[31886] = 8'b11101010;
DRAM[31887] = 8'b11110001;
DRAM[31888] = 8'b11101111;
DRAM[31889] = 8'b11101100;
DRAM[31890] = 8'b11101011;
DRAM[31891] = 8'b11101110;
DRAM[31892] = 8'b11110001;
DRAM[31893] = 8'b11110001;
DRAM[31894] = 8'b11110011;
DRAM[31895] = 8'b11110110;
DRAM[31896] = 8'b11110001;
DRAM[31897] = 8'b11110101;
DRAM[31898] = 8'b11111011;
DRAM[31899] = 8'b11101011;
DRAM[31900] = 8'b11101111;
DRAM[31901] = 8'b11101001;
DRAM[31902] = 8'b11101101;
DRAM[31903] = 8'b11100010;
DRAM[31904] = 8'b11100001;
DRAM[31905] = 8'b11011001;
DRAM[31906] = 8'b11100010;
DRAM[31907] = 8'b11011111;
DRAM[31908] = 8'b11000101;
DRAM[31909] = 8'b10110110;
DRAM[31910] = 8'b10110000;
DRAM[31911] = 8'b10011110;
DRAM[31912] = 8'b10001001;
DRAM[31913] = 8'b10000100;
DRAM[31914] = 8'b10001001;
DRAM[31915] = 8'b1110110;
DRAM[31916] = 8'b1110111;
DRAM[31917] = 8'b10000001;
DRAM[31918] = 8'b1111110;
DRAM[31919] = 8'b1111111;
DRAM[31920] = 8'b10001010;
DRAM[31921] = 8'b10000110;
DRAM[31922] = 8'b10001001;
DRAM[31923] = 8'b10010110;
DRAM[31924] = 8'b10011101;
DRAM[31925] = 8'b10011011;
DRAM[31926] = 8'b10011010;
DRAM[31927] = 8'b10011111;
DRAM[31928] = 8'b10100101;
DRAM[31929] = 8'b10101000;
DRAM[31930] = 8'b10101000;
DRAM[31931] = 8'b10100100;
DRAM[31932] = 8'b10100010;
DRAM[31933] = 8'b10100001;
DRAM[31934] = 8'b10011100;
DRAM[31935] = 8'b10010101;
DRAM[31936] = 8'b10011000;
DRAM[31937] = 8'b10001100;
DRAM[31938] = 8'b10000111;
DRAM[31939] = 8'b1111111;
DRAM[31940] = 8'b1101101;
DRAM[31941] = 8'b1101000;
DRAM[31942] = 8'b1110000;
DRAM[31943] = 8'b1110010;
DRAM[31944] = 8'b1111011;
DRAM[31945] = 8'b10000000;
DRAM[31946] = 8'b10100001;
DRAM[31947] = 8'b11001100;
DRAM[31948] = 8'b11100100;
DRAM[31949] = 8'b11100111;
DRAM[31950] = 8'b11001101;
DRAM[31951] = 8'b10100101;
DRAM[31952] = 8'b1111010;
DRAM[31953] = 8'b10010101;
DRAM[31954] = 8'b10100111;
DRAM[31955] = 8'b10101110;
DRAM[31956] = 8'b11010000;
DRAM[31957] = 8'b11100010;
DRAM[31958] = 8'b11100110;
DRAM[31959] = 8'b11110001;
DRAM[31960] = 8'b11110000;
DRAM[31961] = 8'b11100100;
DRAM[31962] = 8'b10111111;
DRAM[31963] = 8'b10011011;
DRAM[31964] = 8'b10001001;
DRAM[31965] = 8'b10000100;
DRAM[31966] = 8'b10000111;
DRAM[31967] = 8'b10000101;
DRAM[31968] = 8'b10000001;
DRAM[31969] = 8'b10000001;
DRAM[31970] = 8'b10000001;
DRAM[31971] = 8'b10000000;
DRAM[31972] = 8'b10000000;
DRAM[31973] = 8'b10000000;
DRAM[31974] = 8'b1111111;
DRAM[31975] = 8'b1111111;
DRAM[31976] = 8'b1111101;
DRAM[31977] = 8'b1111101;
DRAM[31978] = 8'b1111011;
DRAM[31979] = 8'b1111010;
DRAM[31980] = 8'b1111010;
DRAM[31981] = 8'b1111010;
DRAM[31982] = 8'b1111011;
DRAM[31983] = 8'b1111011;
DRAM[31984] = 8'b1111101;
DRAM[31985] = 8'b1111101;
DRAM[31986] = 8'b1111101;
DRAM[31987] = 8'b1111100;
DRAM[31988] = 8'b1111100;
DRAM[31989] = 8'b1111100;
DRAM[31990] = 8'b1111011;
DRAM[31991] = 8'b1111011;
DRAM[31992] = 8'b1111000;
DRAM[31993] = 8'b1110111;
DRAM[31994] = 8'b1110111;
DRAM[31995] = 8'b1110110;
DRAM[31996] = 8'b1110101;
DRAM[31997] = 8'b1110100;
DRAM[31998] = 8'b1110100;
DRAM[31999] = 8'b1110011;
DRAM[32000] = 8'b10001100;
DRAM[32001] = 8'b10001100;
DRAM[32002] = 8'b10001100;
DRAM[32003] = 8'b10001100;
DRAM[32004] = 8'b10001100;
DRAM[32005] = 8'b10001100;
DRAM[32006] = 8'b10001100;
DRAM[32007] = 8'b10001100;
DRAM[32008] = 8'b10001100;
DRAM[32009] = 8'b10001101;
DRAM[32010] = 8'b10001110;
DRAM[32011] = 8'b10001111;
DRAM[32012] = 8'b10001111;
DRAM[32013] = 8'b10001111;
DRAM[32014] = 8'b10001111;
DRAM[32015] = 8'b10001110;
DRAM[32016] = 8'b10001111;
DRAM[32017] = 8'b10001111;
DRAM[32018] = 8'b10001111;
DRAM[32019] = 8'b10001111;
DRAM[32020] = 8'b10001111;
DRAM[32021] = 8'b10010000;
DRAM[32022] = 8'b10010001;
DRAM[32023] = 8'b10010001;
DRAM[32024] = 8'b10010010;
DRAM[32025] = 8'b10010010;
DRAM[32026] = 8'b10010010;
DRAM[32027] = 8'b10010011;
DRAM[32028] = 8'b10010011;
DRAM[32029] = 8'b10010011;
DRAM[32030] = 8'b10010100;
DRAM[32031] = 8'b10010100;
DRAM[32032] = 8'b10010100;
DRAM[32033] = 8'b10010100;
DRAM[32034] = 8'b10010100;
DRAM[32035] = 8'b10010101;
DRAM[32036] = 8'b10010101;
DRAM[32037] = 8'b10010101;
DRAM[32038] = 8'b10010101;
DRAM[32039] = 8'b10010101;
DRAM[32040] = 8'b10011001;
DRAM[32041] = 8'b10001101;
DRAM[32042] = 8'b10100001;
DRAM[32043] = 8'b10100010;
DRAM[32044] = 8'b10010111;
DRAM[32045] = 8'b10100111;
DRAM[32046] = 8'b10111001;
DRAM[32047] = 8'b11000111;
DRAM[32048] = 8'b10110000;
DRAM[32049] = 8'b10110100;
DRAM[32050] = 8'b10100010;
DRAM[32051] = 8'b10101010;
DRAM[32052] = 8'b10100000;
DRAM[32053] = 8'b10101000;
DRAM[32054] = 8'b10111101;
DRAM[32055] = 8'b11001100;
DRAM[32056] = 8'b11001000;
DRAM[32057] = 8'b11011011;
DRAM[32058] = 8'b11000111;
DRAM[32059] = 8'b11011110;
DRAM[32060] = 8'b11011010;
DRAM[32061] = 8'b11010010;
DRAM[32062] = 8'b11010001;
DRAM[32063] = 8'b10111000;
DRAM[32064] = 8'b10110001;
DRAM[32065] = 8'b10110011;
DRAM[32066] = 8'b10101001;
DRAM[32067] = 8'b10001111;
DRAM[32068] = 8'b10010100;
DRAM[32069] = 8'b10000110;
DRAM[32070] = 8'b1111011;
DRAM[32071] = 8'b1110000;
DRAM[32072] = 8'b1101111;
DRAM[32073] = 8'b1101100;
DRAM[32074] = 8'b1101110;
DRAM[32075] = 8'b1110011;
DRAM[32076] = 8'b1110110;
DRAM[32077] = 8'b1110101;
DRAM[32078] = 8'b1111000;
DRAM[32079] = 8'b1111100;
DRAM[32080] = 8'b10000010;
DRAM[32081] = 8'b10000110;
DRAM[32082] = 8'b10001101;
DRAM[32083] = 8'b10010101;
DRAM[32084] = 8'b10011011;
DRAM[32085] = 8'b10100001;
DRAM[32086] = 8'b10100110;
DRAM[32087] = 8'b10101010;
DRAM[32088] = 8'b10100000;
DRAM[32089] = 8'b10100001;
DRAM[32090] = 8'b10101000;
DRAM[32091] = 8'b10101000;
DRAM[32092] = 8'b10100100;
DRAM[32093] = 8'b10101110;
DRAM[32094] = 8'b10111001;
DRAM[32095] = 8'b10110110;
DRAM[32096] = 8'b10101010;
DRAM[32097] = 8'b10010111;
DRAM[32098] = 8'b10011100;
DRAM[32099] = 8'b1011111;
DRAM[32100] = 8'b111110;
DRAM[32101] = 8'b1000110;
DRAM[32102] = 8'b101001;
DRAM[32103] = 8'b111001;
DRAM[32104] = 8'b101110;
DRAM[32105] = 8'b101100;
DRAM[32106] = 8'b101000;
DRAM[32107] = 8'b101000;
DRAM[32108] = 8'b101101;
DRAM[32109] = 8'b101111;
DRAM[32110] = 8'b100110;
DRAM[32111] = 8'b11001;
DRAM[32112] = 8'b11100;
DRAM[32113] = 8'b101000;
DRAM[32114] = 8'b100000;
DRAM[32115] = 8'b101111;
DRAM[32116] = 8'b111101;
DRAM[32117] = 8'b111001;
DRAM[32118] = 8'b1010110;
DRAM[32119] = 8'b1111001;
DRAM[32120] = 8'b10000100;
DRAM[32121] = 8'b10011110;
DRAM[32122] = 8'b10110110;
DRAM[32123] = 8'b10111100;
DRAM[32124] = 8'b10110011;
DRAM[32125] = 8'b10101101;
DRAM[32126] = 8'b10110110;
DRAM[32127] = 8'b11000101;
DRAM[32128] = 8'b11001011;
DRAM[32129] = 8'b11010010;
DRAM[32130] = 8'b11011010;
DRAM[32131] = 8'b11100000;
DRAM[32132] = 8'b11100111;
DRAM[32133] = 8'b11101111;
DRAM[32134] = 8'b11110010;
DRAM[32135] = 8'b11110010;
DRAM[32136] = 8'b11101111;
DRAM[32137] = 8'b11110101;
DRAM[32138] = 8'b11101111;
DRAM[32139] = 8'b11101010;
DRAM[32140] = 8'b11101101;
DRAM[32141] = 8'b11101100;
DRAM[32142] = 8'b11101101;
DRAM[32143] = 8'b11111000;
DRAM[32144] = 8'b11110000;
DRAM[32145] = 8'b11101110;
DRAM[32146] = 8'b11101101;
DRAM[32147] = 8'b11101101;
DRAM[32148] = 8'b11101111;
DRAM[32149] = 8'b11110001;
DRAM[32150] = 8'b11110100;
DRAM[32151] = 8'b11110111;
DRAM[32152] = 8'b11110001;
DRAM[32153] = 8'b11111000;
DRAM[32154] = 8'b11111111;
DRAM[32155] = 8'b11101001;
DRAM[32156] = 8'b11110110;
DRAM[32157] = 8'b11110000;
DRAM[32158] = 8'b11110111;
DRAM[32159] = 8'b11100011;
DRAM[32160] = 8'b11100111;
DRAM[32161] = 8'b11011110;
DRAM[32162] = 8'b11100000;
DRAM[32163] = 8'b11100101;
DRAM[32164] = 8'b11011111;
DRAM[32165] = 8'b11010010;
DRAM[32166] = 8'b11000001;
DRAM[32167] = 8'b10101111;
DRAM[32168] = 8'b10010111;
DRAM[32169] = 8'b10001001;
DRAM[32170] = 8'b10010000;
DRAM[32171] = 8'b10000010;
DRAM[32172] = 8'b10010100;
DRAM[32173] = 8'b10010111;
DRAM[32174] = 8'b10000010;
DRAM[32175] = 8'b1101100;
DRAM[32176] = 8'b10000110;
DRAM[32177] = 8'b10001110;
DRAM[32178] = 8'b10010011;
DRAM[32179] = 8'b10010110;
DRAM[32180] = 8'b10011011;
DRAM[32181] = 8'b10011111;
DRAM[32182] = 8'b10010110;
DRAM[32183] = 8'b10001000;
DRAM[32184] = 8'b10100000;
DRAM[32185] = 8'b10100111;
DRAM[32186] = 8'b10101100;
DRAM[32187] = 8'b10101100;
DRAM[32188] = 8'b10101100;
DRAM[32189] = 8'b10101011;
DRAM[32190] = 8'b10100101;
DRAM[32191] = 8'b10011110;
DRAM[32192] = 8'b10011100;
DRAM[32193] = 8'b10001111;
DRAM[32194] = 8'b10001010;
DRAM[32195] = 8'b10000011;
DRAM[32196] = 8'b1110001;
DRAM[32197] = 8'b1101011;
DRAM[32198] = 8'b1110001;
DRAM[32199] = 8'b1110010;
DRAM[32200] = 8'b10010000;
DRAM[32201] = 8'b10010000;
DRAM[32202] = 8'b10101101;
DRAM[32203] = 8'b11010111;
DRAM[32204] = 8'b11101010;
DRAM[32205] = 8'b11100110;
DRAM[32206] = 8'b11010100;
DRAM[32207] = 8'b10111111;
DRAM[32208] = 8'b1111011;
DRAM[32209] = 8'b10000100;
DRAM[32210] = 8'b10011111;
DRAM[32211] = 8'b10100010;
DRAM[32212] = 8'b11000011;
DRAM[32213] = 8'b11011000;
DRAM[32214] = 8'b11100101;
DRAM[32215] = 8'b11110101;
DRAM[32216] = 8'b11101011;
DRAM[32217] = 8'b11101010;
DRAM[32218] = 8'b10111100;
DRAM[32219] = 8'b10010111;
DRAM[32220] = 8'b10001000;
DRAM[32221] = 8'b10000001;
DRAM[32222] = 8'b10000110;
DRAM[32223] = 8'b10000011;
DRAM[32224] = 8'b10000010;
DRAM[32225] = 8'b10000001;
DRAM[32226] = 8'b10000001;
DRAM[32227] = 8'b10000001;
DRAM[32228] = 8'b10000000;
DRAM[32229] = 8'b10000000;
DRAM[32230] = 8'b10000000;
DRAM[32231] = 8'b10000000;
DRAM[32232] = 8'b1111110;
DRAM[32233] = 8'b1111100;
DRAM[32234] = 8'b1111011;
DRAM[32235] = 8'b1111001;
DRAM[32236] = 8'b1111001;
DRAM[32237] = 8'b1111001;
DRAM[32238] = 8'b1111011;
DRAM[32239] = 8'b1111011;
DRAM[32240] = 8'b1111110;
DRAM[32241] = 8'b1111110;
DRAM[32242] = 8'b1111101;
DRAM[32243] = 8'b1111101;
DRAM[32244] = 8'b1111101;
DRAM[32245] = 8'b1111100;
DRAM[32246] = 8'b1111100;
DRAM[32247] = 8'b1111100;
DRAM[32248] = 8'b1110111;
DRAM[32249] = 8'b1110111;
DRAM[32250] = 8'b1110111;
DRAM[32251] = 8'b1110110;
DRAM[32252] = 8'b1110101;
DRAM[32253] = 8'b1110100;
DRAM[32254] = 8'b1110100;
DRAM[32255] = 8'b1110011;
DRAM[32256] = 8'b10001101;
DRAM[32257] = 8'b10001101;
DRAM[32258] = 8'b10001101;
DRAM[32259] = 8'b10001101;
DRAM[32260] = 8'b10001101;
DRAM[32261] = 8'b10001101;
DRAM[32262] = 8'b10001101;
DRAM[32263] = 8'b10001101;
DRAM[32264] = 8'b10001101;
DRAM[32265] = 8'b10001110;
DRAM[32266] = 8'b10001110;
DRAM[32267] = 8'b10001111;
DRAM[32268] = 8'b10010000;
DRAM[32269] = 8'b10010000;
DRAM[32270] = 8'b10001111;
DRAM[32271] = 8'b10001111;
DRAM[32272] = 8'b10010000;
DRAM[32273] = 8'b10001111;
DRAM[32274] = 8'b10001111;
DRAM[32275] = 8'b10001111;
DRAM[32276] = 8'b10001111;
DRAM[32277] = 8'b10010000;
DRAM[32278] = 8'b10010001;
DRAM[32279] = 8'b10010010;
DRAM[32280] = 8'b10010001;
DRAM[32281] = 8'b10010001;
DRAM[32282] = 8'b10010010;
DRAM[32283] = 8'b10010010;
DRAM[32284] = 8'b10010010;
DRAM[32285] = 8'b10010011;
DRAM[32286] = 8'b10010011;
DRAM[32287] = 8'b10010011;
DRAM[32288] = 8'b10010101;
DRAM[32289] = 8'b10010110;
DRAM[32290] = 8'b10010110;
DRAM[32291] = 8'b10010111;
DRAM[32292] = 8'b10010111;
DRAM[32293] = 8'b10011000;
DRAM[32294] = 8'b10011000;
DRAM[32295] = 8'b10011000;
DRAM[32296] = 8'b10011010;
DRAM[32297] = 8'b10010100;
DRAM[32298] = 8'b10100010;
DRAM[32299] = 8'b10011001;
DRAM[32300] = 8'b10011100;
DRAM[32301] = 8'b10110000;
DRAM[32302] = 8'b10110001;
DRAM[32303] = 8'b10111110;
DRAM[32304] = 8'b10110001;
DRAM[32305] = 8'b10111000;
DRAM[32306] = 8'b10100010;
DRAM[32307] = 8'b10101111;
DRAM[32308] = 8'b10100001;
DRAM[32309] = 8'b10101010;
DRAM[32310] = 8'b10111001;
DRAM[32311] = 8'b11000111;
DRAM[32312] = 8'b11001101;
DRAM[32313] = 8'b11010101;
DRAM[32314] = 8'b11001100;
DRAM[32315] = 8'b11011011;
DRAM[32316] = 8'b11010001;
DRAM[32317] = 8'b11010101;
DRAM[32318] = 8'b11000010;
DRAM[32319] = 8'b10110111;
DRAM[32320] = 8'b10101001;
DRAM[32321] = 8'b10101111;
DRAM[32322] = 8'b10101000;
DRAM[32323] = 8'b10001100;
DRAM[32324] = 8'b10011000;
DRAM[32325] = 8'b10000101;
DRAM[32326] = 8'b1111100;
DRAM[32327] = 8'b1110100;
DRAM[32328] = 8'b1110101;
DRAM[32329] = 8'b1110001;
DRAM[32330] = 8'b1110000;
DRAM[32331] = 8'b1110011;
DRAM[32332] = 8'b1110100;
DRAM[32333] = 8'b1110100;
DRAM[32334] = 8'b1110110;
DRAM[32335] = 8'b1111011;
DRAM[32336] = 8'b10000101;
DRAM[32337] = 8'b10000100;
DRAM[32338] = 8'b10000101;
DRAM[32339] = 8'b10001001;
DRAM[32340] = 8'b10010000;
DRAM[32341] = 8'b10011011;
DRAM[32342] = 8'b10100101;
DRAM[32343] = 8'b10101011;
DRAM[32344] = 8'b10100000;
DRAM[32345] = 8'b10100010;
DRAM[32346] = 8'b10101100;
DRAM[32347] = 8'b10110001;
DRAM[32348] = 8'b10101111;
DRAM[32349] = 8'b10111000;
DRAM[32350] = 8'b11000010;
DRAM[32351] = 8'b10111111;
DRAM[32352] = 8'b10110110;
DRAM[32353] = 8'b10100111;
DRAM[32354] = 8'b10100001;
DRAM[32355] = 8'b1111101;
DRAM[32356] = 8'b1100011;
DRAM[32357] = 8'b1010111;
DRAM[32358] = 8'b111101;
DRAM[32359] = 8'b111100;
DRAM[32360] = 8'b101101;
DRAM[32361] = 8'b110100;
DRAM[32362] = 8'b111010;
DRAM[32363] = 8'b111100;
DRAM[32364] = 8'b111100;
DRAM[32365] = 8'b111010;
DRAM[32366] = 8'b110010;
DRAM[32367] = 8'b101000;
DRAM[32368] = 8'b1000010;
DRAM[32369] = 8'b1001011;
DRAM[32370] = 8'b1001010;
DRAM[32371] = 8'b1001111;
DRAM[32372] = 8'b1001010;
DRAM[32373] = 8'b1010000;
DRAM[32374] = 8'b1111001;
DRAM[32375] = 8'b10001100;
DRAM[32376] = 8'b10010001;
DRAM[32377] = 8'b10111010;
DRAM[32378] = 8'b11000110;
DRAM[32379] = 8'b10110110;
DRAM[32380] = 8'b10101110;
DRAM[32381] = 8'b10101111;
DRAM[32382] = 8'b11000001;
DRAM[32383] = 8'b11100000;
DRAM[32384] = 8'b11010011;
DRAM[32385] = 8'b11011110;
DRAM[32386] = 8'b11100101;
DRAM[32387] = 8'b11100101;
DRAM[32388] = 8'b11100111;
DRAM[32389] = 8'b11101111;
DRAM[32390] = 8'b11110111;
DRAM[32391] = 8'b11111010;
DRAM[32392] = 8'b11110010;
DRAM[32393] = 8'b11111000;
DRAM[32394] = 8'b11110100;
DRAM[32395] = 8'b11110000;
DRAM[32396] = 8'b11110011;
DRAM[32397] = 8'b11110001;
DRAM[32398] = 8'b11110001;
DRAM[32399] = 8'b11111001;
DRAM[32400] = 8'b11101111;
DRAM[32401] = 8'b11110000;
DRAM[32402] = 8'b11110000;
DRAM[32403] = 8'b11110000;
DRAM[32404] = 8'b11110000;
DRAM[32405] = 8'b11110010;
DRAM[32406] = 8'b11110100;
DRAM[32407] = 8'b11110101;
DRAM[32408] = 8'b11110101;
DRAM[32409] = 8'b11111000;
DRAM[32410] = 8'b11111001;
DRAM[32411] = 8'b11101111;
DRAM[32412] = 8'b11110001;
DRAM[32413] = 8'b11110010;
DRAM[32414] = 8'b11110010;
DRAM[32415] = 8'b11101001;
DRAM[32416] = 8'b11100101;
DRAM[32417] = 8'b11100001;
DRAM[32418] = 8'b11011100;
DRAM[32419] = 8'b11100010;
DRAM[32420] = 8'b11101100;
DRAM[32421] = 8'b11100010;
DRAM[32422] = 8'b11010000;
DRAM[32423] = 8'b11001011;
DRAM[32424] = 8'b10101110;
DRAM[32425] = 8'b10011111;
DRAM[32426] = 8'b10100001;
DRAM[32427] = 8'b1111111;
DRAM[32428] = 8'b10000111;
DRAM[32429] = 8'b10001110;
DRAM[32430] = 8'b10010111;
DRAM[32431] = 8'b10011001;
DRAM[32432] = 8'b1110100;
DRAM[32433] = 8'b1111110;
DRAM[32434] = 8'b10010000;
DRAM[32435] = 8'b10100001;
DRAM[32436] = 8'b10101010;
DRAM[32437] = 8'b10101000;
DRAM[32438] = 8'b10100000;
DRAM[32439] = 8'b10011010;
DRAM[32440] = 8'b10001110;
DRAM[32441] = 8'b10011001;
DRAM[32442] = 8'b10100011;
DRAM[32443] = 8'b10100111;
DRAM[32444] = 8'b10101000;
DRAM[32445] = 8'b10100110;
DRAM[32446] = 8'b10011111;
DRAM[32447] = 8'b10011000;
DRAM[32448] = 8'b10011001;
DRAM[32449] = 8'b10001110;
DRAM[32450] = 8'b10001010;
DRAM[32451] = 8'b10000101;
DRAM[32452] = 8'b1110100;
DRAM[32453] = 8'b1101101;
DRAM[32454] = 8'b1110001;
DRAM[32455] = 8'b1110000;
DRAM[32456] = 8'b10001110;
DRAM[32457] = 8'b10010011;
DRAM[32458] = 8'b10100110;
DRAM[32459] = 8'b11000111;
DRAM[32460] = 8'b11011110;
DRAM[32461] = 8'b11011011;
DRAM[32462] = 8'b11001000;
DRAM[32463] = 8'b10111010;
DRAM[32464] = 8'b10010101;
DRAM[32465] = 8'b1111111;
DRAM[32466] = 8'b10010111;
DRAM[32467] = 8'b10010101;
DRAM[32468] = 8'b10110011;
DRAM[32469] = 8'b11001011;
DRAM[32470] = 8'b11100010;
DRAM[32471] = 8'b11110000;
DRAM[32472] = 8'b11101001;
DRAM[32473] = 8'b11110010;
DRAM[32474] = 8'b11000000;
DRAM[32475] = 8'b10011001;
DRAM[32476] = 8'b10001101;
DRAM[32477] = 8'b10000010;
DRAM[32478] = 8'b10001000;
DRAM[32479] = 8'b10000010;
DRAM[32480] = 8'b10000010;
DRAM[32481] = 8'b10000010;
DRAM[32482] = 8'b10000001;
DRAM[32483] = 8'b10000001;
DRAM[32484] = 8'b10000001;
DRAM[32485] = 8'b10000000;
DRAM[32486] = 8'b10000000;
DRAM[32487] = 8'b10000000;
DRAM[32488] = 8'b1111111;
DRAM[32489] = 8'b1111110;
DRAM[32490] = 8'b1111011;
DRAM[32491] = 8'b1111010;
DRAM[32492] = 8'b1111001;
DRAM[32493] = 8'b1111010;
DRAM[32494] = 8'b1111100;
DRAM[32495] = 8'b1111101;
DRAM[32496] = 8'b1111101;
DRAM[32497] = 8'b1111100;
DRAM[32498] = 8'b1111100;
DRAM[32499] = 8'b1111100;
DRAM[32500] = 8'b1111011;
DRAM[32501] = 8'b1111011;
DRAM[32502] = 8'b1111011;
DRAM[32503] = 8'b1111010;
DRAM[32504] = 8'b1111001;
DRAM[32505] = 8'b1111000;
DRAM[32506] = 8'b1111000;
DRAM[32507] = 8'b1110111;
DRAM[32508] = 8'b1110110;
DRAM[32509] = 8'b1110101;
DRAM[32510] = 8'b1110101;
DRAM[32511] = 8'b1110101;
DRAM[32512] = 8'b10001101;
DRAM[32513] = 8'b10001101;
DRAM[32514] = 8'b10001101;
DRAM[32515] = 8'b10001101;
DRAM[32516] = 8'b10001101;
DRAM[32517] = 8'b10001101;
DRAM[32518] = 8'b10001101;
DRAM[32519] = 8'b10001101;
DRAM[32520] = 8'b10001101;
DRAM[32521] = 8'b10001110;
DRAM[32522] = 8'b10001111;
DRAM[32523] = 8'b10010000;
DRAM[32524] = 8'b10010000;
DRAM[32525] = 8'b10010000;
DRAM[32526] = 8'b10010000;
DRAM[32527] = 8'b10001111;
DRAM[32528] = 8'b10010000;
DRAM[32529] = 8'b10001111;
DRAM[32530] = 8'b10001111;
DRAM[32531] = 8'b10001111;
DRAM[32532] = 8'b10001111;
DRAM[32533] = 8'b10010000;
DRAM[32534] = 8'b10010001;
DRAM[32535] = 8'b10010010;
DRAM[32536] = 8'b10010000;
DRAM[32537] = 8'b10010000;
DRAM[32538] = 8'b10010000;
DRAM[32539] = 8'b10010001;
DRAM[32540] = 8'b10010001;
DRAM[32541] = 8'b10010010;
DRAM[32542] = 8'b10010010;
DRAM[32543] = 8'b10010010;
DRAM[32544] = 8'b10010110;
DRAM[32545] = 8'b10010110;
DRAM[32546] = 8'b10010111;
DRAM[32547] = 8'b10011000;
DRAM[32548] = 8'b10011001;
DRAM[32549] = 8'b10011010;
DRAM[32550] = 8'b10011010;
DRAM[32551] = 8'b10011011;
DRAM[32552] = 8'b10011001;
DRAM[32553] = 8'b10010111;
DRAM[32554] = 8'b10011111;
DRAM[32555] = 8'b10010000;
DRAM[32556] = 8'b10011100;
DRAM[32557] = 8'b10110001;
DRAM[32558] = 8'b10100011;
DRAM[32559] = 8'b10101011;
DRAM[32560] = 8'b10111101;
DRAM[32561] = 8'b11000010;
DRAM[32562] = 8'b10101010;
DRAM[32563] = 8'b10111001;
DRAM[32564] = 8'b10101000;
DRAM[32565] = 8'b10110000;
DRAM[32566] = 8'b10111000;
DRAM[32567] = 8'b11000010;
DRAM[32568] = 8'b11010101;
DRAM[32569] = 8'b11001111;
DRAM[32570] = 8'b11010101;
DRAM[32571] = 8'b11010110;
DRAM[32572] = 8'b11000111;
DRAM[32573] = 8'b11011000;
DRAM[32574] = 8'b10110010;
DRAM[32575] = 8'b10110111;
DRAM[32576] = 8'b10100001;
DRAM[32577] = 8'b10101011;
DRAM[32578] = 8'b10101000;
DRAM[32579] = 8'b10001011;
DRAM[32580] = 8'b10011100;
DRAM[32581] = 8'b10000111;
DRAM[32582] = 8'b1111110;
DRAM[32583] = 8'b1110111;
DRAM[32584] = 8'b1111000;
DRAM[32585] = 8'b1110011;
DRAM[32586] = 8'b1101111;
DRAM[32587] = 8'b1110001;
DRAM[32588] = 8'b1110010;
DRAM[32589] = 8'b1110010;
DRAM[32590] = 8'b1110111;
DRAM[32591] = 8'b1111101;
DRAM[32592] = 8'b1110111;
DRAM[32593] = 8'b1111011;
DRAM[32594] = 8'b10000011;
DRAM[32595] = 8'b10010000;
DRAM[32596] = 8'b10011011;
DRAM[32597] = 8'b10100001;
DRAM[32598] = 8'b10100000;
DRAM[32599] = 8'b10011101;
DRAM[32600] = 8'b10100110;
DRAM[32601] = 8'b10100101;
DRAM[32602] = 8'b10101101;
DRAM[32603] = 8'b10101110;
DRAM[32604] = 8'b10100101;
DRAM[32605] = 8'b10100101;
DRAM[32606] = 8'b10100111;
DRAM[32607] = 8'b10011111;
DRAM[32608] = 8'b10110000;
DRAM[32609] = 8'b10110011;
DRAM[32610] = 8'b10101101;
DRAM[32611] = 8'b10101101;
DRAM[32612] = 8'b10010111;
DRAM[32613] = 8'b1110100;
DRAM[32614] = 8'b1101000;
DRAM[32615] = 8'b1011111;
DRAM[32616] = 8'b1001010;
DRAM[32617] = 8'b1001101;
DRAM[32618] = 8'b1001001;
DRAM[32619] = 8'b1000000;
DRAM[32620] = 8'b111110;
DRAM[32621] = 8'b1000111;
DRAM[32622] = 8'b1010101;
DRAM[32623] = 8'b1011101;
DRAM[32624] = 8'b1010011;
DRAM[32625] = 8'b1011110;
DRAM[32626] = 8'b1100110;
DRAM[32627] = 8'b1100111;
DRAM[32628] = 8'b1010101;
DRAM[32629] = 8'b1100000;
DRAM[32630] = 8'b10001100;
DRAM[32631] = 8'b10010010;
DRAM[32632] = 8'b10100111;
DRAM[32633] = 8'b11001101;
DRAM[32634] = 8'b11001101;
DRAM[32635] = 8'b11000001;
DRAM[32636] = 8'b11001111;
DRAM[32637] = 8'b11010011;
DRAM[32638] = 8'b11001100;
DRAM[32639] = 8'b11010110;
DRAM[32640] = 8'b11011010;
DRAM[32641] = 8'b11101010;
DRAM[32642] = 8'b11110101;
DRAM[32643] = 8'b11110011;
DRAM[32644] = 8'b11101101;
DRAM[32645] = 8'b11110000;
DRAM[32646] = 8'b11111000;
DRAM[32647] = 8'b11111100;
DRAM[32648] = 8'b11110101;
DRAM[32649] = 8'b11111010;
DRAM[32650] = 8'b11110110;
DRAM[32651] = 8'b11110100;
DRAM[32652] = 8'b11111010;
DRAM[32653] = 8'b11110111;
DRAM[32654] = 8'b11110011;
DRAM[32655] = 8'b11110111;
DRAM[32656] = 8'b11110011;
DRAM[32657] = 8'b11110110;
DRAM[32658] = 8'b11111001;
DRAM[32659] = 8'b11111000;
DRAM[32660] = 8'b11111000;
DRAM[32661] = 8'b11111001;
DRAM[32662] = 8'b11111001;
DRAM[32663] = 8'b11111000;
DRAM[32664] = 8'b11111001;
DRAM[32665] = 8'b11111000;
DRAM[32666] = 8'b11101011;
DRAM[32667] = 8'b11110111;
DRAM[32668] = 8'b11101010;
DRAM[32669] = 8'b11110010;
DRAM[32670] = 8'b11101001;
DRAM[32671] = 8'b11110000;
DRAM[32672] = 8'b11101011;
DRAM[32673] = 8'b11101111;
DRAM[32674] = 8'b11100010;
DRAM[32675] = 8'b11011101;
DRAM[32676] = 8'b11100011;
DRAM[32677] = 8'b11010111;
DRAM[32678] = 8'b11001101;
DRAM[32679] = 8'b11011011;
DRAM[32680] = 8'b10111101;
DRAM[32681] = 8'b10100111;
DRAM[32682] = 8'b10101000;
DRAM[32683] = 8'b10001100;
DRAM[32684] = 8'b10100011;
DRAM[32685] = 8'b10101100;
DRAM[32686] = 8'b10101101;
DRAM[32687] = 8'b10100101;
DRAM[32688] = 8'b10100111;
DRAM[32689] = 8'b10010110;
DRAM[32690] = 8'b10011011;
DRAM[32691] = 8'b10110001;
DRAM[32692] = 8'b10101101;
DRAM[32693] = 8'b10010011;
DRAM[32694] = 8'b10010011;
DRAM[32695] = 8'b10101010;
DRAM[32696] = 8'b10110010;
DRAM[32697] = 8'b10110011;
DRAM[32698] = 8'b10101111;
DRAM[32699] = 8'b10100111;
DRAM[32700] = 8'b10100100;
DRAM[32701] = 8'b10100110;
DRAM[32702] = 8'b10100111;
DRAM[32703] = 8'b10100110;
DRAM[32704] = 8'b10011010;
DRAM[32705] = 8'b10001111;
DRAM[32706] = 8'b10001101;
DRAM[32707] = 8'b10001001;
DRAM[32708] = 8'b1111010;
DRAM[32709] = 8'b1110011;
DRAM[32710] = 8'b1110101;
DRAM[32711] = 8'b1110010;
DRAM[32712] = 8'b10001000;
DRAM[32713] = 8'b10010101;
DRAM[32714] = 8'b10100100;
DRAM[32715] = 8'b11000001;
DRAM[32716] = 8'b11100010;
DRAM[32717] = 8'b11101000;
DRAM[32718] = 8'b11010101;
DRAM[32719] = 8'b11000111;
DRAM[32720] = 8'b10110001;
DRAM[32721] = 8'b10000001;
DRAM[32722] = 8'b10010010;
DRAM[32723] = 8'b10001011;
DRAM[32724] = 8'b10100111;
DRAM[32725] = 8'b11000001;
DRAM[32726] = 8'b11011100;
DRAM[32727] = 8'b11100111;
DRAM[32728] = 8'b11101100;
DRAM[32729] = 8'b11111010;
DRAM[32730] = 8'b11000110;
DRAM[32731] = 8'b10011111;
DRAM[32732] = 8'b10010011;
DRAM[32733] = 8'b10000110;
DRAM[32734] = 8'b10001011;
DRAM[32735] = 8'b10000011;
DRAM[32736] = 8'b10000010;
DRAM[32737] = 8'b10000010;
DRAM[32738] = 8'b10000010;
DRAM[32739] = 8'b10000001;
DRAM[32740] = 8'b10000001;
DRAM[32741] = 8'b10000000;
DRAM[32742] = 8'b10000000;
DRAM[32743] = 8'b10000000;
DRAM[32744] = 8'b10000000;
DRAM[32745] = 8'b1111111;
DRAM[32746] = 8'b1111101;
DRAM[32747] = 8'b1111011;
DRAM[32748] = 8'b1111010;
DRAM[32749] = 8'b1111011;
DRAM[32750] = 8'b1111101;
DRAM[32751] = 8'b1111110;
DRAM[32752] = 8'b1111011;
DRAM[32753] = 8'b1111011;
DRAM[32754] = 8'b1111010;
DRAM[32755] = 8'b1111010;
DRAM[32756] = 8'b1111010;
DRAM[32757] = 8'b1111001;
DRAM[32758] = 8'b1111001;
DRAM[32759] = 8'b1111001;
DRAM[32760] = 8'b1111010;
DRAM[32761] = 8'b1111010;
DRAM[32762] = 8'b1111001;
DRAM[32763] = 8'b1111000;
DRAM[32764] = 8'b1111000;
DRAM[32765] = 8'b1110111;
DRAM[32766] = 8'b1110110;
DRAM[32767] = 8'b1110110;
DRAM[32768] = 8'b10001100;
DRAM[32769] = 8'b10001100;
DRAM[32770] = 8'b10001100;
DRAM[32771] = 8'b10001101;
DRAM[32772] = 8'b10001101;
DRAM[32773] = 8'b10001110;
DRAM[32774] = 8'b10001110;
DRAM[32775] = 8'b10001110;
DRAM[32776] = 8'b10001011;
DRAM[32777] = 8'b10001100;
DRAM[32778] = 8'b10001101;
DRAM[32779] = 8'b10001110;
DRAM[32780] = 8'b10010000;
DRAM[32781] = 8'b10010001;
DRAM[32782] = 8'b10010010;
DRAM[32783] = 8'b10010011;
DRAM[32784] = 8'b10001111;
DRAM[32785] = 8'b10010000;
DRAM[32786] = 8'b10010000;
DRAM[32787] = 8'b10010001;
DRAM[32788] = 8'b10010010;
DRAM[32789] = 8'b10010011;
DRAM[32790] = 8'b10010100;
DRAM[32791] = 8'b10010100;
DRAM[32792] = 8'b10010011;
DRAM[32793] = 8'b10010011;
DRAM[32794] = 8'b10010011;
DRAM[32795] = 8'b10010100;
DRAM[32796] = 8'b10010100;
DRAM[32797] = 8'b10010100;
DRAM[32798] = 8'b10010101;
DRAM[32799] = 8'b10010101;
DRAM[32800] = 8'b10010101;
DRAM[32801] = 8'b10010101;
DRAM[32802] = 8'b10010101;
DRAM[32803] = 8'b10010101;
DRAM[32804] = 8'b10010101;
DRAM[32805] = 8'b10010101;
DRAM[32806] = 8'b10010101;
DRAM[32807] = 8'b10010101;
DRAM[32808] = 8'b10011001;
DRAM[32809] = 8'b10011000;
DRAM[32810] = 8'b10010110;
DRAM[32811] = 8'b10010110;
DRAM[32812] = 8'b10011001;
DRAM[32813] = 8'b10011111;
DRAM[32814] = 8'b10100101;
DRAM[32815] = 8'b10101000;
DRAM[32816] = 8'b10110010;
DRAM[32817] = 8'b10101011;
DRAM[32818] = 8'b11001010;
DRAM[32819] = 8'b10111011;
DRAM[32820] = 8'b10101100;
DRAM[32821] = 8'b10110100;
DRAM[32822] = 8'b10100111;
DRAM[32823] = 8'b11001001;
DRAM[32824] = 8'b11001000;
DRAM[32825] = 8'b11001110;
DRAM[32826] = 8'b10111110;
DRAM[32827] = 8'b11001100;
DRAM[32828] = 8'b11000101;
DRAM[32829] = 8'b11000111;
DRAM[32830] = 8'b10101100;
DRAM[32831] = 8'b10101100;
DRAM[32832] = 8'b10101110;
DRAM[32833] = 8'b10100011;
DRAM[32834] = 8'b10011010;
DRAM[32835] = 8'b10010101;
DRAM[32836] = 8'b10001110;
DRAM[32837] = 8'b10000101;
DRAM[32838] = 8'b10000010;
DRAM[32839] = 8'b10000101;
DRAM[32840] = 8'b1110100;
DRAM[32841] = 8'b1110011;
DRAM[32842] = 8'b1110011;
DRAM[32843] = 8'b1110011;
DRAM[32844] = 8'b1110101;
DRAM[32845] = 8'b1110111;
DRAM[32846] = 8'b1111001;
DRAM[32847] = 8'b1111011;
DRAM[32848] = 8'b10000001;
DRAM[32849] = 8'b10000110;
DRAM[32850] = 8'b10010010;
DRAM[32851] = 8'b10011111;
DRAM[32852] = 8'b10100011;
DRAM[32853] = 8'b10100000;
DRAM[32854] = 8'b10011111;
DRAM[32855] = 8'b10100001;
DRAM[32856] = 8'b10100010;
DRAM[32857] = 8'b10100100;
DRAM[32858] = 8'b10101100;
DRAM[32859] = 8'b10110110;
DRAM[32860] = 8'b10110111;
DRAM[32861] = 8'b10110010;
DRAM[32862] = 8'b10110000;
DRAM[32863] = 8'b10110010;
DRAM[32864] = 8'b10101100;
DRAM[32865] = 8'b10101001;
DRAM[32866] = 8'b10010110;
DRAM[32867] = 8'b10000100;
DRAM[32868] = 8'b10010000;
DRAM[32869] = 8'b10100000;
DRAM[32870] = 8'b10000111;
DRAM[32871] = 8'b1011011;
DRAM[32872] = 8'b1100010;
DRAM[32873] = 8'b1100100;
DRAM[32874] = 8'b1010010;
DRAM[32875] = 8'b1001001;
DRAM[32876] = 8'b1100010;
DRAM[32877] = 8'b1011100;
DRAM[32878] = 8'b1101100;
DRAM[32879] = 8'b1001000;
DRAM[32880] = 8'b1001011;
DRAM[32881] = 8'b1011111;
DRAM[32882] = 8'b1111001;
DRAM[32883] = 8'b1101111;
DRAM[32884] = 8'b1111000;
DRAM[32885] = 8'b1111011;
DRAM[32886] = 8'b10010101;
DRAM[32887] = 8'b10011011;
DRAM[32888] = 8'b10111010;
DRAM[32889] = 8'b11000011;
DRAM[32890] = 8'b11000111;
DRAM[32891] = 8'b11000011;
DRAM[32892] = 8'b11000010;
DRAM[32893] = 8'b11001111;
DRAM[32894] = 8'b11100110;
DRAM[32895] = 8'b11111000;
DRAM[32896] = 8'b11101010;
DRAM[32897] = 8'b11101100;
DRAM[32898] = 8'b11110000;
DRAM[32899] = 8'b11110011;
DRAM[32900] = 8'b11110101;
DRAM[32901] = 8'b11110110;
DRAM[32902] = 8'b11110101;
DRAM[32903] = 8'b11110101;
DRAM[32904] = 8'b11110111;
DRAM[32905] = 8'b11110111;
DRAM[32906] = 8'b11110100;
DRAM[32907] = 8'b11110001;
DRAM[32908] = 8'b11110101;
DRAM[32909] = 8'b11111100;
DRAM[32910] = 8'b11111010;
DRAM[32911] = 8'b11110010;
DRAM[32912] = 8'b11110101;
DRAM[32913] = 8'b11110011;
DRAM[32914] = 8'b11110010;
DRAM[32915] = 8'b11110001;
DRAM[32916] = 8'b11110010;
DRAM[32917] = 8'b11110100;
DRAM[32918] = 8'b11110110;
DRAM[32919] = 8'b11111000;
DRAM[32920] = 8'b11110100;
DRAM[32921] = 8'b11110011;
DRAM[32922] = 8'b11110010;
DRAM[32923] = 8'b11110100;
DRAM[32924] = 8'b11110110;
DRAM[32925] = 8'b11110111;
DRAM[32926] = 8'b11110110;
DRAM[32927] = 8'b11110101;
DRAM[32928] = 8'b11110111;
DRAM[32929] = 8'b11110101;
DRAM[32930] = 8'b11110001;
DRAM[32931] = 8'b11101110;
DRAM[32932] = 8'b11101001;
DRAM[32933] = 8'b11100011;
DRAM[32934] = 8'b11011011;
DRAM[32935] = 8'b11010110;
DRAM[32936] = 8'b11011001;
DRAM[32937] = 8'b10111100;
DRAM[32938] = 8'b10101010;
DRAM[32939] = 8'b10100110;
DRAM[32940] = 8'b10100001;
DRAM[32941] = 8'b10011111;
DRAM[32942] = 8'b10011111;
DRAM[32943] = 8'b10011001;
DRAM[32944] = 8'b10011101;
DRAM[32945] = 8'b10101010;
DRAM[32946] = 8'b10011010;
DRAM[32947] = 8'b10001110;
DRAM[32948] = 8'b10101000;
DRAM[32949] = 8'b10110111;
DRAM[32950] = 8'b10101100;
DRAM[32951] = 8'b10100101;
DRAM[32952] = 8'b10101110;
DRAM[32953] = 8'b10100011;
DRAM[32954] = 8'b10011111;
DRAM[32955] = 8'b10101000;
DRAM[32956] = 8'b10110001;
DRAM[32957] = 8'b10101110;
DRAM[32958] = 8'b10100100;
DRAM[32959] = 8'b10011110;
DRAM[32960] = 8'b10010001;
DRAM[32961] = 8'b10001011;
DRAM[32962] = 8'b10000101;
DRAM[32963] = 8'b1111111;
DRAM[32964] = 8'b1111000;
DRAM[32965] = 8'b1110101;
DRAM[32966] = 8'b1111011;
DRAM[32967] = 8'b10000100;
DRAM[32968] = 8'b10000101;
DRAM[32969] = 8'b10010101;
DRAM[32970] = 8'b10101111;
DRAM[32971] = 8'b11001010;
DRAM[32972] = 8'b11100001;
DRAM[32973] = 8'b11101001;
DRAM[32974] = 8'b11100000;
DRAM[32975] = 8'b11010010;
DRAM[32976] = 8'b10110110;
DRAM[32977] = 8'b10010010;
DRAM[32978] = 8'b1111111;
DRAM[32979] = 8'b10001010;
DRAM[32980] = 8'b10011111;
DRAM[32981] = 8'b10111011;
DRAM[32982] = 8'b11010110;
DRAM[32983] = 8'b11100000;
DRAM[32984] = 8'b11110110;
DRAM[32985] = 8'b11111000;
DRAM[32986] = 8'b11011000;
DRAM[32987] = 8'b10000001;
DRAM[32988] = 8'b10010111;
DRAM[32989] = 8'b10000101;
DRAM[32990] = 8'b10001110;
DRAM[32991] = 8'b10000100;
DRAM[32992] = 8'b1111110;
DRAM[32993] = 8'b10000101;
DRAM[32994] = 8'b10000111;
DRAM[32995] = 8'b10000001;
DRAM[32996] = 8'b1111110;
DRAM[32997] = 8'b10000011;
DRAM[32998] = 8'b10000100;
DRAM[32999] = 8'b10000001;
DRAM[33000] = 8'b1111111;
DRAM[33001] = 8'b1111111;
DRAM[33002] = 8'b1111111;
DRAM[33003] = 8'b1111110;
DRAM[33004] = 8'b1111110;
DRAM[33005] = 8'b1111101;
DRAM[33006] = 8'b1111101;
DRAM[33007] = 8'b1111101;
DRAM[33008] = 8'b1111011;
DRAM[33009] = 8'b1111011;
DRAM[33010] = 8'b1111010;
DRAM[33011] = 8'b1111010;
DRAM[33012] = 8'b1111010;
DRAM[33013] = 8'b1111010;
DRAM[33014] = 8'b1111001;
DRAM[33015] = 8'b1111001;
DRAM[33016] = 8'b1111000;
DRAM[33017] = 8'b1110111;
DRAM[33018] = 8'b1110110;
DRAM[33019] = 8'b1110101;
DRAM[33020] = 8'b1110101;
DRAM[33021] = 8'b1110101;
DRAM[33022] = 8'b1110101;
DRAM[33023] = 8'b1110110;
DRAM[33024] = 8'b10001101;
DRAM[33025] = 8'b10001101;
DRAM[33026] = 8'b10001101;
DRAM[33027] = 8'b10001101;
DRAM[33028] = 8'b10001101;
DRAM[33029] = 8'b10001110;
DRAM[33030] = 8'b10001110;
DRAM[33031] = 8'b10001110;
DRAM[33032] = 8'b10001101;
DRAM[33033] = 8'b10001101;
DRAM[33034] = 8'b10001110;
DRAM[33035] = 8'b10001111;
DRAM[33036] = 8'b10010000;
DRAM[33037] = 8'b10010001;
DRAM[33038] = 8'b10010010;
DRAM[33039] = 8'b10010010;
DRAM[33040] = 8'b10010000;
DRAM[33041] = 8'b10010000;
DRAM[33042] = 8'b10010001;
DRAM[33043] = 8'b10010010;
DRAM[33044] = 8'b10010011;
DRAM[33045] = 8'b10010100;
DRAM[33046] = 8'b10010100;
DRAM[33047] = 8'b10010101;
DRAM[33048] = 8'b10010011;
DRAM[33049] = 8'b10010011;
DRAM[33050] = 8'b10010100;
DRAM[33051] = 8'b10010100;
DRAM[33052] = 8'b10010101;
DRAM[33053] = 8'b10010101;
DRAM[33054] = 8'b10010101;
DRAM[33055] = 8'b10010101;
DRAM[33056] = 8'b10010101;
DRAM[33057] = 8'b10010101;
DRAM[33058] = 8'b10010101;
DRAM[33059] = 8'b10010101;
DRAM[33060] = 8'b10010101;
DRAM[33061] = 8'b10010101;
DRAM[33062] = 8'b10010101;
DRAM[33063] = 8'b10010101;
DRAM[33064] = 8'b10010100;
DRAM[33065] = 8'b10010101;
DRAM[33066] = 8'b10010110;
DRAM[33067] = 8'b10010111;
DRAM[33068] = 8'b10011010;
DRAM[33069] = 8'b10011101;
DRAM[33070] = 8'b10011111;
DRAM[33071] = 8'b10100001;
DRAM[33072] = 8'b10101110;
DRAM[33073] = 8'b10101000;
DRAM[33074] = 8'b11001100;
DRAM[33075] = 8'b10111010;
DRAM[33076] = 8'b10110100;
DRAM[33077] = 8'b10110100;
DRAM[33078] = 8'b10101101;
DRAM[33079] = 8'b11001001;
DRAM[33080] = 8'b11001000;
DRAM[33081] = 8'b11010000;
DRAM[33082] = 8'b11000100;
DRAM[33083] = 8'b11001010;
DRAM[33084] = 8'b10111101;
DRAM[33085] = 8'b10111001;
DRAM[33086] = 8'b10100011;
DRAM[33087] = 8'b10101001;
DRAM[33088] = 8'b10100111;
DRAM[33089] = 8'b10011101;
DRAM[33090] = 8'b10010111;
DRAM[33091] = 8'b10010111;
DRAM[33092] = 8'b10010100;
DRAM[33093] = 8'b10001010;
DRAM[33094] = 8'b10000000;
DRAM[33095] = 8'b1111100;
DRAM[33096] = 8'b1111100;
DRAM[33097] = 8'b1111011;
DRAM[33098] = 8'b1111001;
DRAM[33099] = 8'b1111000;
DRAM[33100] = 8'b1111000;
DRAM[33101] = 8'b1111000;
DRAM[33102] = 8'b1111001;
DRAM[33103] = 8'b1111010;
DRAM[33104] = 8'b1110110;
DRAM[33105] = 8'b1111111;
DRAM[33106] = 8'b10010000;
DRAM[33107] = 8'b10100001;
DRAM[33108] = 8'b10101001;
DRAM[33109] = 8'b10101001;
DRAM[33110] = 8'b10101000;
DRAM[33111] = 8'b10101010;
DRAM[33112] = 8'b10100111;
DRAM[33113] = 8'b10101011;
DRAM[33114] = 8'b10101111;
DRAM[33115] = 8'b10110000;
DRAM[33116] = 8'b10110000;
DRAM[33117] = 8'b10101101;
DRAM[33118] = 8'b10101010;
DRAM[33119] = 8'b10101000;
DRAM[33120] = 8'b10101001;
DRAM[33121] = 8'b10100111;
DRAM[33122] = 8'b10100010;
DRAM[33123] = 8'b10011111;
DRAM[33124] = 8'b10100010;
DRAM[33125] = 8'b10100010;
DRAM[33126] = 8'b10010100;
DRAM[33127] = 8'b10000010;
DRAM[33128] = 8'b10000111;
DRAM[33129] = 8'b1111110;
DRAM[33130] = 8'b1101110;
DRAM[33131] = 8'b1111000;
DRAM[33132] = 8'b1110100;
DRAM[33133] = 8'b1101001;
DRAM[33134] = 8'b1101001;
DRAM[33135] = 8'b1101010;
DRAM[33136] = 8'b1101001;
DRAM[33137] = 8'b1101111;
DRAM[33138] = 8'b1111111;
DRAM[33139] = 8'b1111000;
DRAM[33140] = 8'b10001001;
DRAM[33141] = 8'b10001100;
DRAM[33142] = 8'b10100011;
DRAM[33143] = 8'b10101001;
DRAM[33144] = 8'b11001111;
DRAM[33145] = 8'b11001010;
DRAM[33146] = 8'b11001001;
DRAM[33147] = 8'b11001111;
DRAM[33148] = 8'b11011001;
DRAM[33149] = 8'b11100011;
DRAM[33150] = 8'b11101011;
DRAM[33151] = 8'b11110000;
DRAM[33152] = 8'b11110110;
DRAM[33153] = 8'b11110110;
DRAM[33154] = 8'b11110111;
DRAM[33155] = 8'b11110111;
DRAM[33156] = 8'b11110111;
DRAM[33157] = 8'b11110110;
DRAM[33158] = 8'b11110100;
DRAM[33159] = 8'b11110011;
DRAM[33160] = 8'b11110110;
DRAM[33161] = 8'b11110110;
DRAM[33162] = 8'b11110011;
DRAM[33163] = 8'b11110001;
DRAM[33164] = 8'b11110101;
DRAM[33165] = 8'b11111100;
DRAM[33166] = 8'b11111010;
DRAM[33167] = 8'b11110100;
DRAM[33168] = 8'b11110101;
DRAM[33169] = 8'b11110100;
DRAM[33170] = 8'b11110010;
DRAM[33171] = 8'b11110001;
DRAM[33172] = 8'b11110010;
DRAM[33173] = 8'b11110100;
DRAM[33174] = 8'b11110110;
DRAM[33175] = 8'b11110111;
DRAM[33176] = 8'b11110100;
DRAM[33177] = 8'b11110100;
DRAM[33178] = 8'b11110100;
DRAM[33179] = 8'b11110110;
DRAM[33180] = 8'b11111010;
DRAM[33181] = 8'b11111100;
DRAM[33182] = 8'b11111100;
DRAM[33183] = 8'b11111011;
DRAM[33184] = 8'b11110101;
DRAM[33185] = 8'b11110011;
DRAM[33186] = 8'b11110001;
DRAM[33187] = 8'b11101110;
DRAM[33188] = 8'b11101011;
DRAM[33189] = 8'b11100101;
DRAM[33190] = 8'b11011111;
DRAM[33191] = 8'b11011010;
DRAM[33192] = 8'b11001111;
DRAM[33193] = 8'b11001001;
DRAM[33194] = 8'b11001000;
DRAM[33195] = 8'b10111111;
DRAM[33196] = 8'b10101010;
DRAM[33197] = 8'b10100101;
DRAM[33198] = 8'b10110000;
DRAM[33199] = 8'b10110110;
DRAM[33200] = 8'b10101111;
DRAM[33201] = 8'b10000011;
DRAM[33202] = 8'b10010010;
DRAM[33203] = 8'b10110110;
DRAM[33204] = 8'b10100111;
DRAM[33205] = 8'b10100000;
DRAM[33206] = 8'b10111001;
DRAM[33207] = 8'b11000101;
DRAM[33208] = 8'b10101000;
DRAM[33209] = 8'b10101001;
DRAM[33210] = 8'b10101110;
DRAM[33211] = 8'b10110000;
DRAM[33212] = 8'b10101010;
DRAM[33213] = 8'b10100000;
DRAM[33214] = 8'b10011111;
DRAM[33215] = 8'b10100101;
DRAM[33216] = 8'b10100100;
DRAM[33217] = 8'b10011001;
DRAM[33218] = 8'b10001110;
DRAM[33219] = 8'b10000110;
DRAM[33220] = 8'b10000000;
DRAM[33221] = 8'b1111010;
DRAM[33222] = 8'b1111010;
DRAM[33223] = 8'b1111110;
DRAM[33224] = 8'b10010000;
DRAM[33225] = 8'b10011101;
DRAM[33226] = 8'b10110010;
DRAM[33227] = 8'b11001101;
DRAM[33228] = 8'b11100011;
DRAM[33229] = 8'b11101000;
DRAM[33230] = 8'b11010111;
DRAM[33231] = 8'b11000010;
DRAM[33232] = 8'b10010100;
DRAM[33233] = 8'b10010010;
DRAM[33234] = 8'b10001110;
DRAM[33235] = 8'b10000010;
DRAM[33236] = 8'b10000100;
DRAM[33237] = 8'b10100101;
DRAM[33238] = 8'b11000111;
DRAM[33239] = 8'b11001101;
DRAM[33240] = 8'b11011010;
DRAM[33241] = 8'b11110100;
DRAM[33242] = 8'b11011001;
DRAM[33243] = 8'b10010011;
DRAM[33244] = 8'b10001111;
DRAM[33245] = 8'b10001100;
DRAM[33246] = 8'b10001011;
DRAM[33247] = 8'b10000111;
DRAM[33248] = 8'b10000101;
DRAM[33249] = 8'b10000001;
DRAM[33250] = 8'b1111101;
DRAM[33251] = 8'b1111101;
DRAM[33252] = 8'b10000010;
DRAM[33253] = 8'b10000110;
DRAM[33254] = 8'b10000001;
DRAM[33255] = 8'b1111010;
DRAM[33256] = 8'b1111111;
DRAM[33257] = 8'b1111111;
DRAM[33258] = 8'b1111111;
DRAM[33259] = 8'b1111110;
DRAM[33260] = 8'b1111110;
DRAM[33261] = 8'b1111110;
DRAM[33262] = 8'b1111101;
DRAM[33263] = 8'b1111101;
DRAM[33264] = 8'b1111011;
DRAM[33265] = 8'b1111011;
DRAM[33266] = 8'b1111011;
DRAM[33267] = 8'b1111010;
DRAM[33268] = 8'b1111010;
DRAM[33269] = 8'b1111010;
DRAM[33270] = 8'b1111001;
DRAM[33271] = 8'b1111001;
DRAM[33272] = 8'b1111000;
DRAM[33273] = 8'b1110111;
DRAM[33274] = 8'b1110110;
DRAM[33275] = 8'b1110110;
DRAM[33276] = 8'b1110101;
DRAM[33277] = 8'b1110101;
DRAM[33278] = 8'b1110110;
DRAM[33279] = 8'b1110110;
DRAM[33280] = 8'b10001110;
DRAM[33281] = 8'b10001110;
DRAM[33282] = 8'b10001110;
DRAM[33283] = 8'b10001110;
DRAM[33284] = 8'b10001110;
DRAM[33285] = 8'b10001110;
DRAM[33286] = 8'b10001101;
DRAM[33287] = 8'b10001101;
DRAM[33288] = 8'b10001111;
DRAM[33289] = 8'b10001111;
DRAM[33290] = 8'b10001111;
DRAM[33291] = 8'b10010000;
DRAM[33292] = 8'b10010001;
DRAM[33293] = 8'b10010001;
DRAM[33294] = 8'b10010001;
DRAM[33295] = 8'b10010010;
DRAM[33296] = 8'b10010001;
DRAM[33297] = 8'b10010010;
DRAM[33298] = 8'b10010010;
DRAM[33299] = 8'b10010011;
DRAM[33300] = 8'b10010100;
DRAM[33301] = 8'b10010100;
DRAM[33302] = 8'b10010101;
DRAM[33303] = 8'b10010101;
DRAM[33304] = 8'b10010100;
DRAM[33305] = 8'b10010100;
DRAM[33306] = 8'b10010101;
DRAM[33307] = 8'b10010101;
DRAM[33308] = 8'b10010101;
DRAM[33309] = 8'b10010110;
DRAM[33310] = 8'b10010110;
DRAM[33311] = 8'b10010110;
DRAM[33312] = 8'b10010110;
DRAM[33313] = 8'b10010110;
DRAM[33314] = 8'b10010110;
DRAM[33315] = 8'b10010110;
DRAM[33316] = 8'b10010110;
DRAM[33317] = 8'b10010110;
DRAM[33318] = 8'b10010110;
DRAM[33319] = 8'b10010110;
DRAM[33320] = 8'b10010010;
DRAM[33321] = 8'b10010100;
DRAM[33322] = 8'b10010111;
DRAM[33323] = 8'b10011010;
DRAM[33324] = 8'b10011100;
DRAM[33325] = 8'b10011100;
DRAM[33326] = 8'b10011011;
DRAM[33327] = 8'b10011011;
DRAM[33328] = 8'b10100011;
DRAM[33329] = 8'b10011100;
DRAM[33330] = 8'b11000110;
DRAM[33331] = 8'b10110001;
DRAM[33332] = 8'b10111011;
DRAM[33333] = 8'b10110001;
DRAM[33334] = 8'b10110001;
DRAM[33335] = 8'b10111111;
DRAM[33336] = 8'b11000101;
DRAM[33337] = 8'b11001111;
DRAM[33338] = 8'b11000110;
DRAM[33339] = 8'b11000101;
DRAM[33340] = 8'b10110011;
DRAM[33341] = 8'b10101000;
DRAM[33342] = 8'b10011011;
DRAM[33343] = 8'b10101000;
DRAM[33344] = 8'b10100011;
DRAM[33345] = 8'b10011010;
DRAM[33346] = 8'b10010100;
DRAM[33347] = 8'b10010110;
DRAM[33348] = 8'b10011000;
DRAM[33349] = 8'b10010001;
DRAM[33350] = 8'b10000101;
DRAM[33351] = 8'b1111101;
DRAM[33352] = 8'b10000010;
DRAM[33353] = 8'b10000000;
DRAM[33354] = 8'b1111110;
DRAM[33355] = 8'b1111100;
DRAM[33356] = 8'b1111011;
DRAM[33357] = 8'b1111011;
DRAM[33358] = 8'b1111011;
DRAM[33359] = 8'b1111100;
DRAM[33360] = 8'b1111011;
DRAM[33361] = 8'b10000000;
DRAM[33362] = 8'b10001100;
DRAM[33363] = 8'b10011010;
DRAM[33364] = 8'b10100000;
DRAM[33365] = 8'b10011110;
DRAM[33366] = 8'b10011111;
DRAM[33367] = 8'b10100010;
DRAM[33368] = 8'b10101111;
DRAM[33369] = 8'b10110110;
DRAM[33370] = 8'b10111000;
DRAM[33371] = 8'b10110010;
DRAM[33372] = 8'b10110001;
DRAM[33373] = 8'b10110011;
DRAM[33374] = 8'b10101111;
DRAM[33375] = 8'b10100111;
DRAM[33376] = 8'b10101010;
DRAM[33377] = 8'b10100111;
DRAM[33378] = 8'b10101011;
DRAM[33379] = 8'b10110001;
DRAM[33380] = 8'b10100110;
DRAM[33381] = 8'b10010010;
DRAM[33382] = 8'b10001011;
DRAM[33383] = 8'b10010011;
DRAM[33384] = 8'b10001111;
DRAM[33385] = 8'b10000000;
DRAM[33386] = 8'b1110101;
DRAM[33387] = 8'b10000110;
DRAM[33388] = 8'b1111001;
DRAM[33389] = 8'b10000000;
DRAM[33390] = 8'b1100110;
DRAM[33391] = 8'b1110000;
DRAM[33392] = 8'b10000100;
DRAM[33393] = 8'b1111010;
DRAM[33394] = 8'b10000010;
DRAM[33395] = 8'b10000100;
DRAM[33396] = 8'b10011111;
DRAM[33397] = 8'b10100110;
DRAM[33398] = 8'b10111011;
DRAM[33399] = 8'b11000001;
DRAM[33400] = 8'b11001111;
DRAM[33401] = 8'b11001001;
DRAM[33402] = 8'b11001011;
DRAM[33403] = 8'b11011011;
DRAM[33404] = 8'b11101000;
DRAM[33405] = 8'b11101101;
DRAM[33406] = 8'b11101111;
DRAM[33407] = 8'b11110010;
DRAM[33408] = 8'b11101111;
DRAM[33409] = 8'b11110000;
DRAM[33410] = 8'b11110000;
DRAM[33411] = 8'b11110001;
DRAM[33412] = 8'b11110011;
DRAM[33413] = 8'b11110101;
DRAM[33414] = 8'b11110110;
DRAM[33415] = 8'b11110111;
DRAM[33416] = 8'b11110101;
DRAM[33417] = 8'b11110101;
DRAM[33418] = 8'b11110011;
DRAM[33419] = 8'b11110010;
DRAM[33420] = 8'b11110110;
DRAM[33421] = 8'b11111011;
DRAM[33422] = 8'b11111010;
DRAM[33423] = 8'b11110110;
DRAM[33424] = 8'b11110110;
DRAM[33425] = 8'b11110101;
DRAM[33426] = 8'b11110100;
DRAM[33427] = 8'b11110011;
DRAM[33428] = 8'b11110100;
DRAM[33429] = 8'b11110101;
DRAM[33430] = 8'b11110111;
DRAM[33431] = 8'b11111000;
DRAM[33432] = 8'b11110111;
DRAM[33433] = 8'b11110110;
DRAM[33434] = 8'b11110110;
DRAM[33435] = 8'b11111000;
DRAM[33436] = 8'b11111011;
DRAM[33437] = 8'b11111101;
DRAM[33438] = 8'b11111101;
DRAM[33439] = 8'b11111100;
DRAM[33440] = 8'b11110100;
DRAM[33441] = 8'b11110010;
DRAM[33442] = 8'b11110000;
DRAM[33443] = 8'b11101111;
DRAM[33444] = 8'b11101100;
DRAM[33445] = 8'b11101000;
DRAM[33446] = 8'b11100010;
DRAM[33447] = 8'b11011110;
DRAM[33448] = 8'b11101001;
DRAM[33449] = 8'b11010101;
DRAM[33450] = 8'b11000101;
DRAM[33451] = 8'b10111011;
DRAM[33452] = 8'b10110010;
DRAM[33453] = 8'b10101110;
DRAM[33454] = 8'b10100001;
DRAM[33455] = 8'b10001010;
DRAM[33456] = 8'b11000000;
DRAM[33457] = 8'b10110001;
DRAM[33458] = 8'b10100001;
DRAM[33459] = 8'b10101001;
DRAM[33460] = 8'b10111101;
DRAM[33461] = 8'b10111110;
DRAM[33462] = 8'b10110000;
DRAM[33463] = 8'b10101001;
DRAM[33464] = 8'b10100100;
DRAM[33465] = 8'b10100111;
DRAM[33466] = 8'b10101100;
DRAM[33467] = 8'b10101101;
DRAM[33468] = 8'b10100101;
DRAM[33469] = 8'b10011101;
DRAM[33470] = 8'b10011100;
DRAM[33471] = 8'b10100001;
DRAM[33472] = 8'b10011011;
DRAM[33473] = 8'b10010000;
DRAM[33474] = 8'b10000101;
DRAM[33475] = 8'b10000011;
DRAM[33476] = 8'b10000011;
DRAM[33477] = 8'b10000001;
DRAM[33478] = 8'b10000000;
DRAM[33479] = 8'b10000001;
DRAM[33480] = 8'b10011001;
DRAM[33481] = 8'b10100100;
DRAM[33482] = 8'b10111000;
DRAM[33483] = 8'b11010001;
DRAM[33484] = 8'b11100110;
DRAM[33485] = 8'b11100110;
DRAM[33486] = 8'b11001101;
DRAM[33487] = 8'b10110011;
DRAM[33488] = 8'b10011010;
DRAM[33489] = 8'b10011110;
DRAM[33490] = 8'b10100000;
DRAM[33491] = 8'b10010100;
DRAM[33492] = 8'b10001101;
DRAM[33493] = 8'b10100110;
DRAM[33494] = 8'b11000101;
DRAM[33495] = 8'b11001110;
DRAM[33496] = 8'b11010000;
DRAM[33497] = 8'b11110010;
DRAM[33498] = 8'b11010010;
DRAM[33499] = 8'b10011010;
DRAM[33500] = 8'b1111011;
DRAM[33501] = 8'b10000101;
DRAM[33502] = 8'b10000010;
DRAM[33503] = 8'b10001010;
DRAM[33504] = 8'b10000111;
DRAM[33505] = 8'b10000000;
DRAM[33506] = 8'b1111101;
DRAM[33507] = 8'b10000000;
DRAM[33508] = 8'b10000100;
DRAM[33509] = 8'b10000011;
DRAM[33510] = 8'b1111111;
DRAM[33511] = 8'b1111101;
DRAM[33512] = 8'b1111111;
DRAM[33513] = 8'b1111111;
DRAM[33514] = 8'b1111111;
DRAM[33515] = 8'b1111111;
DRAM[33516] = 8'b1111110;
DRAM[33517] = 8'b1111110;
DRAM[33518] = 8'b1111110;
DRAM[33519] = 8'b1111101;
DRAM[33520] = 8'b1111100;
DRAM[33521] = 8'b1111011;
DRAM[33522] = 8'b1111011;
DRAM[33523] = 8'b1111011;
DRAM[33524] = 8'b1111010;
DRAM[33525] = 8'b1111010;
DRAM[33526] = 8'b1111001;
DRAM[33527] = 8'b1111001;
DRAM[33528] = 8'b1111000;
DRAM[33529] = 8'b1111000;
DRAM[33530] = 8'b1110111;
DRAM[33531] = 8'b1110110;
DRAM[33532] = 8'b1110101;
DRAM[33533] = 8'b1110101;
DRAM[33534] = 8'b1110110;
DRAM[33535] = 8'b1110110;
DRAM[33536] = 8'b10001111;
DRAM[33537] = 8'b10001111;
DRAM[33538] = 8'b10001111;
DRAM[33539] = 8'b10001111;
DRAM[33540] = 8'b10001110;
DRAM[33541] = 8'b10001110;
DRAM[33542] = 8'b10001110;
DRAM[33543] = 8'b10001110;
DRAM[33544] = 8'b10010001;
DRAM[33545] = 8'b10010001;
DRAM[33546] = 8'b10010001;
DRAM[33547] = 8'b10010001;
DRAM[33548] = 8'b10010001;
DRAM[33549] = 8'b10010010;
DRAM[33550] = 8'b10010010;
DRAM[33551] = 8'b10010010;
DRAM[33552] = 8'b10010011;
DRAM[33553] = 8'b10010011;
DRAM[33554] = 8'b10010100;
DRAM[33555] = 8'b10010100;
DRAM[33556] = 8'b10010101;
DRAM[33557] = 8'b10010101;
DRAM[33558] = 8'b10010110;
DRAM[33559] = 8'b10010110;
DRAM[33560] = 8'b10010101;
DRAM[33561] = 8'b10010101;
DRAM[33562] = 8'b10010110;
DRAM[33563] = 8'b10010110;
DRAM[33564] = 8'b10010111;
DRAM[33565] = 8'b10010111;
DRAM[33566] = 8'b10010111;
DRAM[33567] = 8'b10010111;
DRAM[33568] = 8'b10010111;
DRAM[33569] = 8'b10010111;
DRAM[33570] = 8'b10010111;
DRAM[33571] = 8'b10010111;
DRAM[33572] = 8'b10010111;
DRAM[33573] = 8'b10010111;
DRAM[33574] = 8'b10010111;
DRAM[33575] = 8'b10010111;
DRAM[33576] = 8'b10010110;
DRAM[33577] = 8'b10011000;
DRAM[33578] = 8'b10011011;
DRAM[33579] = 8'b10011101;
DRAM[33580] = 8'b10011101;
DRAM[33581] = 8'b10011101;
DRAM[33582] = 8'b10011100;
DRAM[33583] = 8'b10011011;
DRAM[33584] = 8'b10011111;
DRAM[33585] = 8'b10010101;
DRAM[33586] = 8'b10111011;
DRAM[33587] = 8'b10100111;
DRAM[33588] = 8'b11000011;
DRAM[33589] = 8'b10110101;
DRAM[33590] = 8'b10111000;
DRAM[33591] = 8'b10110111;
DRAM[33592] = 8'b11000011;
DRAM[33593] = 8'b11001001;
DRAM[33594] = 8'b11000010;
DRAM[33595] = 8'b10111101;
DRAM[33596] = 8'b10101111;
DRAM[33597] = 8'b10011111;
DRAM[33598] = 8'b10011001;
DRAM[33599] = 8'b10101001;
DRAM[33600] = 8'b10011111;
DRAM[33601] = 8'b10011010;
DRAM[33602] = 8'b10010101;
DRAM[33603] = 8'b10010110;
DRAM[33604] = 8'b10010111;
DRAM[33605] = 8'b10010100;
DRAM[33606] = 8'b10001110;
DRAM[33607] = 8'b10001001;
DRAM[33608] = 8'b10000001;
DRAM[33609] = 8'b10000000;
DRAM[33610] = 8'b1111110;
DRAM[33611] = 8'b1111100;
DRAM[33612] = 8'b1111100;
DRAM[33613] = 8'b1111101;
DRAM[33614] = 8'b1111110;
DRAM[33615] = 8'b1111110;
DRAM[33616] = 8'b10000011;
DRAM[33617] = 8'b10000100;
DRAM[33618] = 8'b10001001;
DRAM[33619] = 8'b10010000;
DRAM[33620] = 8'b10010100;
DRAM[33621] = 8'b10010100;
DRAM[33622] = 8'b10010111;
DRAM[33623] = 8'b10011101;
DRAM[33624] = 8'b10100010;
DRAM[33625] = 8'b10101110;
DRAM[33626] = 8'b10110000;
DRAM[33627] = 8'b10101001;
DRAM[33628] = 8'b10101010;
DRAM[33629] = 8'b10110001;
DRAM[33630] = 8'b10101100;
DRAM[33631] = 8'b10011110;
DRAM[33632] = 8'b10100111;
DRAM[33633] = 8'b10100011;
DRAM[33634] = 8'b10100111;
DRAM[33635] = 8'b10101100;
DRAM[33636] = 8'b10100000;
DRAM[33637] = 8'b10001010;
DRAM[33638] = 8'b10000111;
DRAM[33639] = 8'b10010011;
DRAM[33640] = 8'b10010000;
DRAM[33641] = 8'b10001111;
DRAM[33642] = 8'b10010111;
DRAM[33643] = 8'b10001011;
DRAM[33644] = 8'b1111110;
DRAM[33645] = 8'b10010001;
DRAM[33646] = 8'b1111000;
DRAM[33647] = 8'b1111101;
DRAM[33648] = 8'b10010100;
DRAM[33649] = 8'b10000100;
DRAM[33650] = 8'b10001011;
DRAM[33651] = 8'b10010010;
DRAM[33652] = 8'b10110000;
DRAM[33653] = 8'b10110010;
DRAM[33654] = 8'b11000101;
DRAM[33655] = 8'b11001010;
DRAM[33656] = 8'b11001101;
DRAM[33657] = 8'b11001110;
DRAM[33658] = 8'b11011000;
DRAM[33659] = 8'b11100111;
DRAM[33660] = 8'b11101010;
DRAM[33661] = 8'b11100101;
DRAM[33662] = 8'b11101011;
DRAM[33663] = 8'b11110111;
DRAM[33664] = 8'b11101100;
DRAM[33665] = 8'b11101100;
DRAM[33666] = 8'b11101100;
DRAM[33667] = 8'b11101101;
DRAM[33668] = 8'b11110000;
DRAM[33669] = 8'b11110011;
DRAM[33670] = 8'b11110111;
DRAM[33671] = 8'b11111001;
DRAM[33672] = 8'b11110110;
DRAM[33673] = 8'b11110101;
DRAM[33674] = 8'b11110100;
DRAM[33675] = 8'b11110100;
DRAM[33676] = 8'b11110111;
DRAM[33677] = 8'b11111011;
DRAM[33678] = 8'b11111011;
DRAM[33679] = 8'b11111001;
DRAM[33680] = 8'b11111001;
DRAM[33681] = 8'b11111001;
DRAM[33682] = 8'b11111000;
DRAM[33683] = 8'b11110111;
DRAM[33684] = 8'b11110111;
DRAM[33685] = 8'b11111000;
DRAM[33686] = 8'b11111001;
DRAM[33687] = 8'b11111010;
DRAM[33688] = 8'b11111011;
DRAM[33689] = 8'b11111010;
DRAM[33690] = 8'b11111000;
DRAM[33691] = 8'b11111000;
DRAM[33692] = 8'b11111001;
DRAM[33693] = 8'b11111001;
DRAM[33694] = 8'b11111000;
DRAM[33695] = 8'b11110110;
DRAM[33696] = 8'b11110100;
DRAM[33697] = 8'b11110010;
DRAM[33698] = 8'b11110001;
DRAM[33699] = 8'b11101111;
DRAM[33700] = 8'b11101101;
DRAM[33701] = 8'b11101001;
DRAM[33702] = 8'b11100100;
DRAM[33703] = 8'b11011111;
DRAM[33704] = 8'b11011010;
DRAM[33705] = 8'b11011101;
DRAM[33706] = 8'b11100001;
DRAM[33707] = 8'b11010100;
DRAM[33708] = 8'b10111101;
DRAM[33709] = 8'b10110110;
DRAM[33710] = 8'b10110100;
DRAM[33711] = 8'b10101010;
DRAM[33712] = 8'b1101110;
DRAM[33713] = 8'b10101001;
DRAM[33714] = 8'b10101110;
DRAM[33715] = 8'b10010100;
DRAM[33716] = 8'b10100001;
DRAM[33717] = 8'b10101111;
DRAM[33718] = 8'b10100111;
DRAM[33719] = 8'b10100110;
DRAM[33720] = 8'b10101011;
DRAM[33721] = 8'b10100011;
DRAM[33722] = 8'b10011111;
DRAM[33723] = 8'b10100100;
DRAM[33724] = 8'b10101101;
DRAM[33725] = 8'b10101101;
DRAM[33726] = 8'b10100011;
DRAM[33727] = 8'b10011001;
DRAM[33728] = 8'b10001010;
DRAM[33729] = 8'b10000010;
DRAM[33730] = 8'b1111101;
DRAM[33731] = 8'b1111110;
DRAM[33732] = 8'b10000010;
DRAM[33733] = 8'b10000100;
DRAM[33734] = 8'b10000111;
DRAM[33735] = 8'b10001100;
DRAM[33736] = 8'b10011011;
DRAM[33737] = 8'b10101001;
DRAM[33738] = 8'b11000000;
DRAM[33739] = 8'b11011000;
DRAM[33740] = 8'b11101000;
DRAM[33741] = 8'b11100011;
DRAM[33742] = 8'b11001001;
DRAM[33743] = 8'b10101111;
DRAM[33744] = 8'b10100101;
DRAM[33745] = 8'b10001110;
DRAM[33746] = 8'b10001010;
DRAM[33747] = 8'b10010111;
DRAM[33748] = 8'b10011011;
DRAM[33749] = 8'b10100100;
DRAM[33750] = 8'b10111010;
DRAM[33751] = 8'b11001010;
DRAM[33752] = 8'b11011000;
DRAM[33753] = 8'b11101011;
DRAM[33754] = 8'b11010000;
DRAM[33755] = 8'b10100111;
DRAM[33756] = 8'b10000111;
DRAM[33757] = 8'b10000100;
DRAM[33758] = 8'b1111101;
DRAM[33759] = 8'b10000100;
DRAM[33760] = 8'b10000010;
DRAM[33761] = 8'b10000001;
DRAM[33762] = 8'b10000100;
DRAM[33763] = 8'b10000111;
DRAM[33764] = 8'b10000011;
DRAM[33765] = 8'b1111101;
DRAM[33766] = 8'b1111111;
DRAM[33767] = 8'b10001000;
DRAM[33768] = 8'b10000000;
DRAM[33769] = 8'b10000000;
DRAM[33770] = 8'b1111111;
DRAM[33771] = 8'b1111111;
DRAM[33772] = 8'b1111111;
DRAM[33773] = 8'b1111110;
DRAM[33774] = 8'b1111110;
DRAM[33775] = 8'b1111110;
DRAM[33776] = 8'b1111101;
DRAM[33777] = 8'b1111100;
DRAM[33778] = 8'b1111100;
DRAM[33779] = 8'b1111011;
DRAM[33780] = 8'b1111010;
DRAM[33781] = 8'b1111010;
DRAM[33782] = 8'b1111001;
DRAM[33783] = 8'b1111001;
DRAM[33784] = 8'b1111001;
DRAM[33785] = 8'b1111000;
DRAM[33786] = 8'b1110111;
DRAM[33787] = 8'b1110110;
DRAM[33788] = 8'b1110110;
DRAM[33789] = 8'b1110110;
DRAM[33790] = 8'b1110110;
DRAM[33791] = 8'b1110111;
DRAM[33792] = 8'b10010000;
DRAM[33793] = 8'b10010000;
DRAM[33794] = 8'b10010000;
DRAM[33795] = 8'b10001111;
DRAM[33796] = 8'b10001111;
DRAM[33797] = 8'b10001111;
DRAM[33798] = 8'b10001111;
DRAM[33799] = 8'b10001111;
DRAM[33800] = 8'b10010010;
DRAM[33801] = 8'b10010010;
DRAM[33802] = 8'b10010010;
DRAM[33803] = 8'b10010011;
DRAM[33804] = 8'b10010011;
DRAM[33805] = 8'b10010011;
DRAM[33806] = 8'b10010011;
DRAM[33807] = 8'b10010011;
DRAM[33808] = 8'b10010101;
DRAM[33809] = 8'b10010101;
DRAM[33810] = 8'b10010101;
DRAM[33811] = 8'b10010101;
DRAM[33812] = 8'b10010110;
DRAM[33813] = 8'b10010110;
DRAM[33814] = 8'b10010110;
DRAM[33815] = 8'b10010110;
DRAM[33816] = 8'b10010111;
DRAM[33817] = 8'b10010111;
DRAM[33818] = 8'b10010111;
DRAM[33819] = 8'b10010111;
DRAM[33820] = 8'b10011000;
DRAM[33821] = 8'b10011000;
DRAM[33822] = 8'b10011001;
DRAM[33823] = 8'b10011001;
DRAM[33824] = 8'b10011001;
DRAM[33825] = 8'b10011001;
DRAM[33826] = 8'b10011001;
DRAM[33827] = 8'b10011001;
DRAM[33828] = 8'b10011001;
DRAM[33829] = 8'b10011001;
DRAM[33830] = 8'b10011001;
DRAM[33831] = 8'b10011001;
DRAM[33832] = 8'b10011011;
DRAM[33833] = 8'b10011011;
DRAM[33834] = 8'b10011010;
DRAM[33835] = 8'b10011010;
DRAM[33836] = 8'b10011011;
DRAM[33837] = 8'b10011100;
DRAM[33838] = 8'b10011100;
DRAM[33839] = 8'b10011101;
DRAM[33840] = 8'b10100101;
DRAM[33841] = 8'b10011000;
DRAM[33842] = 8'b10110011;
DRAM[33843] = 8'b10100101;
DRAM[33844] = 8'b11001001;
DRAM[33845] = 8'b10111110;
DRAM[33846] = 8'b11000011;
DRAM[33847] = 8'b10110110;
DRAM[33848] = 8'b11000111;
DRAM[33849] = 8'b11000100;
DRAM[33850] = 8'b10111101;
DRAM[33851] = 8'b10110100;
DRAM[33852] = 8'b10101111;
DRAM[33853] = 8'b10011011;
DRAM[33854] = 8'b10010111;
DRAM[33855] = 8'b10100100;
DRAM[33856] = 8'b10010101;
DRAM[33857] = 8'b10011001;
DRAM[33858] = 8'b10011101;
DRAM[33859] = 8'b10011100;
DRAM[33860] = 8'b10011001;
DRAM[33861] = 8'b10010101;
DRAM[33862] = 8'b10010001;
DRAM[33863] = 8'b10001110;
DRAM[33864] = 8'b10000001;
DRAM[33865] = 8'b10000000;
DRAM[33866] = 8'b1111110;
DRAM[33867] = 8'b1111011;
DRAM[33868] = 8'b1111010;
DRAM[33869] = 8'b1111010;
DRAM[33870] = 8'b1111010;
DRAM[33871] = 8'b1111011;
DRAM[33872] = 8'b1111000;
DRAM[33873] = 8'b1111100;
DRAM[33874] = 8'b10000111;
DRAM[33875] = 8'b10010011;
DRAM[33876] = 8'b10011010;
DRAM[33877] = 8'b10011100;
DRAM[33878] = 8'b10100000;
DRAM[33879] = 8'b10100110;
DRAM[33880] = 8'b10100011;
DRAM[33881] = 8'b10101111;
DRAM[33882] = 8'b10110011;
DRAM[33883] = 8'b10101110;
DRAM[33884] = 8'b10110000;
DRAM[33885] = 8'b10110110;
DRAM[33886] = 8'b10101111;
DRAM[33887] = 8'b10100000;
DRAM[33888] = 8'b10011111;
DRAM[33889] = 8'b10011101;
DRAM[33890] = 8'b10011100;
DRAM[33891] = 8'b10011111;
DRAM[33892] = 8'b10100000;
DRAM[33893] = 8'b10011101;
DRAM[33894] = 8'b10011101;
DRAM[33895] = 8'b10011110;
DRAM[33896] = 8'b10011011;
DRAM[33897] = 8'b10010111;
DRAM[33898] = 8'b10101011;
DRAM[33899] = 8'b10000101;
DRAM[33900] = 8'b1111010;
DRAM[33901] = 8'b1111011;
DRAM[33902] = 8'b1111101;
DRAM[33903] = 8'b10001110;
DRAM[33904] = 8'b10011100;
DRAM[33905] = 8'b10010010;
DRAM[33906] = 8'b10011101;
DRAM[33907] = 8'b10100011;
DRAM[33908] = 8'b10111011;
DRAM[33909] = 8'b10110101;
DRAM[33910] = 8'b11000011;
DRAM[33911] = 8'b11000111;
DRAM[33912] = 8'b11011001;
DRAM[33913] = 8'b11011010;
DRAM[33914] = 8'b11100001;
DRAM[33915] = 8'b11101001;
DRAM[33916] = 8'b11101001;
DRAM[33917] = 8'b11100100;
DRAM[33918] = 8'b11100111;
DRAM[33919] = 8'b11110000;
DRAM[33920] = 8'b11111010;
DRAM[33921] = 8'b11111001;
DRAM[33922] = 8'b11110110;
DRAM[33923] = 8'b11110100;
DRAM[33924] = 8'b11110100;
DRAM[33925] = 8'b11110101;
DRAM[33926] = 8'b11111000;
DRAM[33927] = 8'b11111001;
DRAM[33928] = 8'b11111000;
DRAM[33929] = 8'b11110110;
DRAM[33930] = 8'b11110110;
DRAM[33931] = 8'b11110111;
DRAM[33932] = 8'b11111001;
DRAM[33933] = 8'b11111010;
DRAM[33934] = 8'b11111011;
DRAM[33935] = 8'b11111100;
DRAM[33936] = 8'b11111101;
DRAM[33937] = 8'b11111100;
DRAM[33938] = 8'b11111100;
DRAM[33939] = 8'b11111011;
DRAM[33940] = 8'b11111011;
DRAM[33941] = 8'b11111100;
DRAM[33942] = 8'b11111100;
DRAM[33943] = 8'b11111100;
DRAM[33944] = 8'b11111100;
DRAM[33945] = 8'b11111010;
DRAM[33946] = 8'b11111001;
DRAM[33947] = 8'b11111001;
DRAM[33948] = 8'b11111010;
DRAM[33949] = 8'b11111010;
DRAM[33950] = 8'b11111001;
DRAM[33951] = 8'b11110111;
DRAM[33952] = 8'b11110110;
DRAM[33953] = 8'b11110100;
DRAM[33954] = 8'b11110011;
DRAM[33955] = 8'b11110001;
DRAM[33956] = 8'b11101111;
DRAM[33957] = 8'b11101010;
DRAM[33958] = 8'b11100100;
DRAM[33959] = 8'b11100000;
DRAM[33960] = 8'b11011010;
DRAM[33961] = 8'b11011110;
DRAM[33962] = 8'b11100110;
DRAM[33963] = 8'b11100000;
DRAM[33964] = 8'b11001110;
DRAM[33965] = 8'b11000111;
DRAM[33966] = 8'b11000110;
DRAM[33967] = 8'b10111110;
DRAM[33968] = 8'b10110000;
DRAM[33969] = 8'b10100111;
DRAM[33970] = 8'b10111010;
DRAM[33971] = 8'b11000000;
DRAM[33972] = 8'b10100011;
DRAM[33973] = 8'b10011110;
DRAM[33974] = 8'b10100111;
DRAM[33975] = 8'b10010111;
DRAM[33976] = 8'b10110010;
DRAM[33977] = 8'b10101000;
DRAM[33978] = 8'b10100000;
DRAM[33979] = 8'b10100101;
DRAM[33980] = 8'b10110010;
DRAM[33981] = 8'b10110110;
DRAM[33982] = 8'b10101000;
DRAM[33983] = 8'b10011000;
DRAM[33984] = 8'b10001100;
DRAM[33985] = 8'b10001000;
DRAM[33986] = 8'b10000101;
DRAM[33987] = 8'b10000100;
DRAM[33988] = 8'b10000010;
DRAM[33989] = 8'b10000010;
DRAM[33990] = 8'b10001001;
DRAM[33991] = 8'b10010010;
DRAM[33992] = 8'b10011101;
DRAM[33993] = 8'b10110000;
DRAM[33994] = 8'b11001011;
DRAM[33995] = 8'b11011111;
DRAM[33996] = 8'b11101000;
DRAM[33997] = 8'b11100000;
DRAM[33998] = 8'b11001001;
DRAM[33999] = 8'b10110011;
DRAM[34000] = 8'b10011110;
DRAM[34001] = 8'b10000010;
DRAM[34002] = 8'b1111100;
DRAM[34003] = 8'b10001111;
DRAM[34004] = 8'b10011011;
DRAM[34005] = 8'b10100111;
DRAM[34006] = 8'b10111100;
DRAM[34007] = 8'b11001011;
DRAM[34008] = 8'b11011011;
DRAM[34009] = 8'b11010100;
DRAM[34010] = 8'b11001010;
DRAM[34011] = 8'b10110100;
DRAM[34012] = 8'b10101100;
DRAM[34013] = 8'b10010011;
DRAM[34014] = 8'b10001001;
DRAM[34015] = 8'b10000101;
DRAM[34016] = 8'b10000011;
DRAM[34017] = 8'b10000001;
DRAM[34018] = 8'b10000010;
DRAM[34019] = 8'b10000101;
DRAM[34020] = 8'b10000100;
DRAM[34021] = 8'b10000001;
DRAM[34022] = 8'b10000010;
DRAM[34023] = 8'b10000101;
DRAM[34024] = 8'b10000000;
DRAM[34025] = 8'b10000000;
DRAM[34026] = 8'b10000000;
DRAM[34027] = 8'b1111111;
DRAM[34028] = 8'b1111111;
DRAM[34029] = 8'b1111111;
DRAM[34030] = 8'b1111110;
DRAM[34031] = 8'b1111110;
DRAM[34032] = 8'b1111110;
DRAM[34033] = 8'b1111101;
DRAM[34034] = 8'b1111101;
DRAM[34035] = 8'b1111100;
DRAM[34036] = 8'b1111011;
DRAM[34037] = 8'b1111010;
DRAM[34038] = 8'b1111001;
DRAM[34039] = 8'b1111001;
DRAM[34040] = 8'b1111001;
DRAM[34041] = 8'b1111000;
DRAM[34042] = 8'b1110111;
DRAM[34043] = 8'b1110111;
DRAM[34044] = 8'b1110110;
DRAM[34045] = 8'b1110110;
DRAM[34046] = 8'b1110111;
DRAM[34047] = 8'b1110111;
DRAM[34048] = 8'b10001111;
DRAM[34049] = 8'b10001111;
DRAM[34050] = 8'b10001111;
DRAM[34051] = 8'b10010000;
DRAM[34052] = 8'b10010000;
DRAM[34053] = 8'b10010001;
DRAM[34054] = 8'b10010001;
DRAM[34055] = 8'b10010001;
DRAM[34056] = 8'b10010010;
DRAM[34057] = 8'b10010011;
DRAM[34058] = 8'b10010011;
DRAM[34059] = 8'b10010011;
DRAM[34060] = 8'b10010100;
DRAM[34061] = 8'b10010101;
DRAM[34062] = 8'b10010101;
DRAM[34063] = 8'b10010101;
DRAM[34064] = 8'b10010111;
DRAM[34065] = 8'b10010111;
DRAM[34066] = 8'b10010111;
DRAM[34067] = 8'b10010111;
DRAM[34068] = 8'b10010111;
DRAM[34069] = 8'b10010111;
DRAM[34070] = 8'b10010111;
DRAM[34071] = 8'b10010111;
DRAM[34072] = 8'b10011000;
DRAM[34073] = 8'b10011000;
DRAM[34074] = 8'b10011000;
DRAM[34075] = 8'b10011001;
DRAM[34076] = 8'b10011001;
DRAM[34077] = 8'b10011001;
DRAM[34078] = 8'b10011010;
DRAM[34079] = 8'b10011010;
DRAM[34080] = 8'b10011010;
DRAM[34081] = 8'b10011010;
DRAM[34082] = 8'b10011010;
DRAM[34083] = 8'b10011010;
DRAM[34084] = 8'b10011010;
DRAM[34085] = 8'b10011010;
DRAM[34086] = 8'b10011010;
DRAM[34087] = 8'b10011010;
DRAM[34088] = 8'b10011100;
DRAM[34089] = 8'b10011010;
DRAM[34090] = 8'b10011000;
DRAM[34091] = 8'b10010111;
DRAM[34092] = 8'b10011000;
DRAM[34093] = 8'b10011001;
DRAM[34094] = 8'b10011100;
DRAM[34095] = 8'b10011101;
DRAM[34096] = 8'b10100011;
DRAM[34097] = 8'b10011011;
DRAM[34098] = 8'b10101000;
DRAM[34099] = 8'b10100001;
DRAM[34100] = 8'b11000000;
DRAM[34101] = 8'b10111100;
DRAM[34102] = 8'b11000100;
DRAM[34103] = 8'b10110110;
DRAM[34104] = 8'b11001011;
DRAM[34105] = 8'b11000001;
DRAM[34106] = 8'b10111011;
DRAM[34107] = 8'b10101110;
DRAM[34108] = 8'b10110000;
DRAM[34109] = 8'b10010101;
DRAM[34110] = 8'b10010011;
DRAM[34111] = 8'b10011101;
DRAM[34112] = 8'b10010000;
DRAM[34113] = 8'b10011100;
DRAM[34114] = 8'b10100110;
DRAM[34115] = 8'b10100101;
DRAM[34116] = 8'b10011111;
DRAM[34117] = 8'b10011000;
DRAM[34118] = 8'b10010000;
DRAM[34119] = 8'b10001010;
DRAM[34120] = 8'b10000111;
DRAM[34121] = 8'b10000100;
DRAM[34122] = 8'b10000000;
DRAM[34123] = 8'b1111100;
DRAM[34124] = 8'b1111000;
DRAM[34125] = 8'b1110110;
DRAM[34126] = 8'b1110101;
DRAM[34127] = 8'b1110100;
DRAM[34128] = 8'b1101100;
DRAM[34129] = 8'b1110101;
DRAM[34130] = 8'b10001000;
DRAM[34131] = 8'b10011100;
DRAM[34132] = 8'b10100101;
DRAM[34133] = 8'b10100100;
DRAM[34134] = 8'b10100010;
DRAM[34135] = 8'b10100011;
DRAM[34136] = 8'b10101101;
DRAM[34137] = 8'b10110011;
DRAM[34138] = 8'b10110101;
DRAM[34139] = 8'b10110011;
DRAM[34140] = 8'b10110101;
DRAM[34141] = 8'b10110111;
DRAM[34142] = 8'b10101111;
DRAM[34143] = 8'b10100010;
DRAM[34144] = 8'b10100000;
DRAM[34145] = 8'b10011110;
DRAM[34146] = 8'b10011010;
DRAM[34147] = 8'b10011001;
DRAM[34148] = 8'b10100001;
DRAM[34149] = 8'b10101010;
DRAM[34150] = 8'b10101001;
DRAM[34151] = 8'b10100010;
DRAM[34152] = 8'b10101011;
DRAM[34153] = 8'b10000100;
DRAM[34154] = 8'b10000001;
DRAM[34155] = 8'b1110011;
DRAM[34156] = 8'b10000101;
DRAM[34157] = 8'b1110111;
DRAM[34158] = 8'b10000101;
DRAM[34159] = 8'b10010110;
DRAM[34160] = 8'b10010011;
DRAM[34161] = 8'b10010101;
DRAM[34162] = 8'b10101011;
DRAM[34163] = 8'b10110001;
DRAM[34164] = 8'b11000110;
DRAM[34165] = 8'b11000000;
DRAM[34166] = 8'b11001100;
DRAM[34167] = 8'b11001101;
DRAM[34168] = 8'b11010101;
DRAM[34169] = 8'b11010011;
DRAM[34170] = 8'b11010100;
DRAM[34171] = 8'b11011100;
DRAM[34172] = 8'b11100111;
DRAM[34173] = 8'b11101101;
DRAM[34174] = 8'b11101101;
DRAM[34175] = 8'b11101010;
DRAM[34176] = 8'b11111011;
DRAM[34177] = 8'b11111010;
DRAM[34178] = 8'b11111000;
DRAM[34179] = 8'b11111000;
DRAM[34180] = 8'b11111001;
DRAM[34181] = 8'b11111011;
DRAM[34182] = 8'b11111110;
DRAM[34183] = 8'b11111111;
DRAM[34184] = 8'b11111100;
DRAM[34185] = 8'b11111001;
DRAM[34186] = 8'b11111001;
DRAM[34187] = 8'b11111011;
DRAM[34188] = 8'b11111100;
DRAM[34189] = 8'b11111010;
DRAM[34190] = 8'b11111011;
DRAM[34191] = 8'b11111110;
DRAM[34192] = 8'b11111110;
DRAM[34193] = 8'b11111110;
DRAM[34194] = 8'b11111110;
DRAM[34195] = 8'b11111110;
DRAM[34196] = 8'b11111110;
DRAM[34197] = 8'b11111101;
DRAM[34198] = 8'b11111101;
DRAM[34199] = 8'b11111101;
DRAM[34200] = 8'b11111010;
DRAM[34201] = 8'b11111001;
DRAM[34202] = 8'b11111001;
DRAM[34203] = 8'b11111010;
DRAM[34204] = 8'b11111101;
DRAM[34205] = 8'b11111111;
DRAM[34206] = 8'b11111111;
DRAM[34207] = 8'b11111110;
DRAM[34208] = 8'b11111001;
DRAM[34209] = 8'b11110111;
DRAM[34210] = 8'b11110110;
DRAM[34211] = 8'b11110100;
DRAM[34212] = 8'b11110010;
DRAM[34213] = 8'b11101110;
DRAM[34214] = 8'b11101001;
DRAM[34215] = 8'b11100100;
DRAM[34216] = 8'b11101000;
DRAM[34217] = 8'b11010101;
DRAM[34218] = 8'b11010000;
DRAM[34219] = 8'b11010110;
DRAM[34220] = 8'b11010110;
DRAM[34221] = 8'b11010001;
DRAM[34222] = 8'b11000101;
DRAM[34223] = 8'b10110011;
DRAM[34224] = 8'b10111111;
DRAM[34225] = 8'b10010101;
DRAM[34226] = 8'b10000101;
DRAM[34227] = 8'b10011110;
DRAM[34228] = 8'b10110101;
DRAM[34229] = 8'b10110111;
DRAM[34230] = 8'b10101111;
DRAM[34231] = 8'b10100111;
DRAM[34232] = 8'b10101011;
DRAM[34233] = 8'b10101100;
DRAM[34234] = 8'b10101010;
DRAM[34235] = 8'b10101000;
DRAM[34236] = 8'b10101001;
DRAM[34237] = 8'b10101000;
DRAM[34238] = 8'b10100001;
DRAM[34239] = 8'b10011001;
DRAM[34240] = 8'b10001110;
DRAM[34241] = 8'b10001010;
DRAM[34242] = 8'b10001000;
DRAM[34243] = 8'b10000110;
DRAM[34244] = 8'b10000011;
DRAM[34245] = 8'b10000011;
DRAM[34246] = 8'b10001101;
DRAM[34247] = 8'b10011001;
DRAM[34248] = 8'b10100010;
DRAM[34249] = 8'b10110111;
DRAM[34250] = 8'b11010010;
DRAM[34251] = 8'b11100100;
DRAM[34252] = 8'b11101001;
DRAM[34253] = 8'b11100001;
DRAM[34254] = 8'b11001100;
DRAM[34255] = 8'b10111001;
DRAM[34256] = 8'b10010001;
DRAM[34257] = 8'b10001011;
DRAM[34258] = 8'b10001100;
DRAM[34259] = 8'b10001100;
DRAM[34260] = 8'b10010001;
DRAM[34261] = 8'b10101010;
DRAM[34262] = 8'b11000100;
DRAM[34263] = 8'b11001010;
DRAM[34264] = 8'b11001111;
DRAM[34265] = 8'b10111000;
DRAM[34266] = 8'b10101011;
DRAM[34267] = 8'b10011111;
DRAM[34268] = 8'b10100011;
DRAM[34269] = 8'b10011000;
DRAM[34270] = 8'b10011010;
DRAM[34271] = 8'b10010110;
DRAM[34272] = 8'b10001011;
DRAM[34273] = 8'b10000101;
DRAM[34274] = 8'b1111101;
DRAM[34275] = 8'b1111101;
DRAM[34276] = 8'b10000110;
DRAM[34277] = 8'b10001100;
DRAM[34278] = 8'b10000100;
DRAM[34279] = 8'b1111001;
DRAM[34280] = 8'b10000001;
DRAM[34281] = 8'b10000000;
DRAM[34282] = 8'b10000000;
DRAM[34283] = 8'b10000000;
DRAM[34284] = 8'b1111111;
DRAM[34285] = 8'b1111111;
DRAM[34286] = 8'b1111111;
DRAM[34287] = 8'b1111111;
DRAM[34288] = 8'b1111110;
DRAM[34289] = 8'b1111110;
DRAM[34290] = 8'b1111101;
DRAM[34291] = 8'b1111100;
DRAM[34292] = 8'b1111011;
DRAM[34293] = 8'b1111010;
DRAM[34294] = 8'b1111001;
DRAM[34295] = 8'b1111001;
DRAM[34296] = 8'b1111001;
DRAM[34297] = 8'b1111001;
DRAM[34298] = 8'b1111000;
DRAM[34299] = 8'b1110111;
DRAM[34300] = 8'b1110111;
DRAM[34301] = 8'b1110111;
DRAM[34302] = 8'b1110111;
DRAM[34303] = 8'b1110111;
DRAM[34304] = 8'b10001110;
DRAM[34305] = 8'b10001110;
DRAM[34306] = 8'b10001111;
DRAM[34307] = 8'b10010000;
DRAM[34308] = 8'b10010001;
DRAM[34309] = 8'b10010010;
DRAM[34310] = 8'b10010011;
DRAM[34311] = 8'b10010100;
DRAM[34312] = 8'b10010010;
DRAM[34313] = 8'b10010010;
DRAM[34314] = 8'b10010011;
DRAM[34315] = 8'b10010100;
DRAM[34316] = 8'b10010101;
DRAM[34317] = 8'b10010110;
DRAM[34318] = 8'b10010111;
DRAM[34319] = 8'b10010111;
DRAM[34320] = 8'b10011000;
DRAM[34321] = 8'b10011000;
DRAM[34322] = 8'b10011000;
DRAM[34323] = 8'b10011000;
DRAM[34324] = 8'b10011000;
DRAM[34325] = 8'b10011000;
DRAM[34326] = 8'b10011000;
DRAM[34327] = 8'b10010111;
DRAM[34328] = 8'b10011001;
DRAM[34329] = 8'b10011001;
DRAM[34330] = 8'b10011001;
DRAM[34331] = 8'b10011001;
DRAM[34332] = 8'b10011010;
DRAM[34333] = 8'b10011010;
DRAM[34334] = 8'b10011011;
DRAM[34335] = 8'b10011011;
DRAM[34336] = 8'b10011011;
DRAM[34337] = 8'b10011011;
DRAM[34338] = 8'b10011011;
DRAM[34339] = 8'b10011011;
DRAM[34340] = 8'b10011011;
DRAM[34341] = 8'b10011011;
DRAM[34342] = 8'b10011011;
DRAM[34343] = 8'b10011011;
DRAM[34344] = 8'b10011100;
DRAM[34345] = 8'b10011011;
DRAM[34346] = 8'b10011010;
DRAM[34347] = 8'b10011001;
DRAM[34348] = 8'b10011001;
DRAM[34349] = 8'b10011011;
DRAM[34350] = 8'b10011101;
DRAM[34351] = 8'b10011111;
DRAM[34352] = 8'b10011101;
DRAM[34353] = 8'b10100000;
DRAM[34354] = 8'b10100001;
DRAM[34355] = 8'b10011111;
DRAM[34356] = 8'b10101101;
DRAM[34357] = 8'b10110011;
DRAM[34358] = 8'b10111111;
DRAM[34359] = 8'b10111010;
DRAM[34360] = 8'b11000110;
DRAM[34361] = 8'b10111011;
DRAM[34362] = 8'b10111001;
DRAM[34363] = 8'b10101010;
DRAM[34364] = 8'b10101111;
DRAM[34365] = 8'b10001111;
DRAM[34366] = 8'b10010001;
DRAM[34367] = 8'b10011101;
DRAM[34368] = 8'b10100010;
DRAM[34369] = 8'b10101001;
DRAM[34370] = 8'b10101100;
DRAM[34371] = 8'b10100110;
DRAM[34372] = 8'b10100000;
DRAM[34373] = 8'b10011011;
DRAM[34374] = 8'b10010100;
DRAM[34375] = 8'b10001100;
DRAM[34376] = 8'b10001010;
DRAM[34377] = 8'b10001000;
DRAM[34378] = 8'b10000011;
DRAM[34379] = 8'b1111110;
DRAM[34380] = 8'b1111010;
DRAM[34381] = 8'b1110111;
DRAM[34382] = 8'b1110101;
DRAM[34383] = 8'b1110100;
DRAM[34384] = 8'b1110000;
DRAM[34385] = 8'b1111001;
DRAM[34386] = 8'b10001011;
DRAM[34387] = 8'b10011101;
DRAM[34388] = 8'b10100110;
DRAM[34389] = 8'b10100101;
DRAM[34390] = 8'b10100100;
DRAM[34391] = 8'b10100101;
DRAM[34392] = 8'b10101010;
DRAM[34393] = 8'b10101000;
DRAM[34394] = 8'b10100110;
DRAM[34395] = 8'b10100111;
DRAM[34396] = 8'b10101001;
DRAM[34397] = 8'b10101000;
DRAM[34398] = 8'b10100010;
DRAM[34399] = 8'b10011100;
DRAM[34400] = 8'b10100100;
DRAM[34401] = 8'b10100010;
DRAM[34402] = 8'b10011111;
DRAM[34403] = 8'b10100000;
DRAM[34404] = 8'b10100011;
DRAM[34405] = 8'b10100101;
DRAM[34406] = 8'b10100100;
DRAM[34407] = 8'b10100010;
DRAM[34408] = 8'b10101001;
DRAM[34409] = 8'b10001100;
DRAM[34410] = 8'b1111000;
DRAM[34411] = 8'b10001011;
DRAM[34412] = 8'b10011110;
DRAM[34413] = 8'b10010110;
DRAM[34414] = 8'b10100000;
DRAM[34415] = 8'b10100101;
DRAM[34416] = 8'b10001101;
DRAM[34417] = 8'b10011001;
DRAM[34418] = 8'b10110100;
DRAM[34419] = 8'b10111000;
DRAM[34420] = 8'b11001101;
DRAM[34421] = 8'b11001011;
DRAM[34422] = 8'b11010101;
DRAM[34423] = 8'b11001111;
DRAM[34424] = 8'b11000110;
DRAM[34425] = 8'b11001110;
DRAM[34426] = 8'b11010011;
DRAM[34427] = 8'b11010101;
DRAM[34428] = 8'b11100000;
DRAM[34429] = 8'b11101110;
DRAM[34430] = 8'b11110000;
DRAM[34431] = 8'b11101010;
DRAM[34432] = 8'b11110011;
DRAM[34433] = 8'b11110100;
DRAM[34434] = 8'b11110100;
DRAM[34435] = 8'b11110110;
DRAM[34436] = 8'b11111001;
DRAM[34437] = 8'b11111101;
DRAM[34438] = 8'b11111111;
DRAM[34439] = 8'b11111111;
DRAM[34440] = 8'b11111111;
DRAM[34441] = 8'b11111100;
DRAM[34442] = 8'b11111100;
DRAM[34443] = 8'b11111111;
DRAM[34444] = 8'b11111110;
DRAM[34445] = 8'b11111010;
DRAM[34446] = 8'b11111011;
DRAM[34447] = 8'b11111111;
DRAM[34448] = 8'b11111110;
DRAM[34449] = 8'b11111110;
DRAM[34450] = 8'b11111110;
DRAM[34451] = 8'b11111110;
DRAM[34452] = 8'b11111101;
DRAM[34453] = 8'b11111101;
DRAM[34454] = 8'b11111100;
DRAM[34455] = 8'b11111011;
DRAM[34456] = 8'b11111000;
DRAM[34457] = 8'b11110111;
DRAM[34458] = 8'b11110111;
DRAM[34459] = 8'b11111010;
DRAM[34460] = 8'b11111101;
DRAM[34461] = 8'b11111111;
DRAM[34462] = 8'b11111111;
DRAM[34463] = 8'b11111111;
DRAM[34464] = 8'b11111011;
DRAM[34465] = 8'b11111010;
DRAM[34466] = 8'b11111001;
DRAM[34467] = 8'b11111001;
DRAM[34468] = 8'b11111000;
DRAM[34469] = 8'b11110101;
DRAM[34470] = 8'b11110000;
DRAM[34471] = 8'b11101100;
DRAM[34472] = 8'b11011001;
DRAM[34473] = 8'b11010010;
DRAM[34474] = 8'b11011101;
DRAM[34475] = 8'b11100101;
DRAM[34476] = 8'b11010110;
DRAM[34477] = 8'b11001010;
DRAM[34478] = 8'b11010011;
DRAM[34479] = 8'b11011110;
DRAM[34480] = 8'b11001100;
DRAM[34481] = 8'b11010010;
DRAM[34482] = 8'b10110100;
DRAM[34483] = 8'b10100100;
DRAM[34484] = 8'b10110100;
DRAM[34485] = 8'b10101001;
DRAM[34486] = 8'b10011110;
DRAM[34487] = 8'b10111000;
DRAM[34488] = 8'b10100101;
DRAM[34489] = 8'b10101100;
DRAM[34490] = 8'b10101111;
DRAM[34491] = 8'b10101001;
DRAM[34492] = 8'b10100100;
DRAM[34493] = 8'b10100010;
DRAM[34494] = 8'b10011111;
DRAM[34495] = 8'b10011011;
DRAM[34496] = 8'b10001111;
DRAM[34497] = 8'b10001000;
DRAM[34498] = 8'b10000011;
DRAM[34499] = 8'b10000010;
DRAM[34500] = 8'b10000100;
DRAM[34501] = 8'b10001000;
DRAM[34502] = 8'b10010010;
DRAM[34503] = 8'b10011100;
DRAM[34504] = 8'b10100101;
DRAM[34505] = 8'b10110111;
DRAM[34506] = 8'b11010000;
DRAM[34507] = 8'b11100011;
DRAM[34508] = 8'b11101110;
DRAM[34509] = 8'b11101001;
DRAM[34510] = 8'b11010110;
DRAM[34511] = 8'b11000100;
DRAM[34512] = 8'b10010100;
DRAM[34513] = 8'b10001100;
DRAM[34514] = 8'b10001010;
DRAM[34515] = 8'b10000111;
DRAM[34516] = 8'b10000100;
DRAM[34517] = 8'b10010100;
DRAM[34518] = 8'b10100111;
DRAM[34519] = 8'b10101011;
DRAM[34520] = 8'b10101011;
DRAM[34521] = 8'b10100011;
DRAM[34522] = 8'b10001111;
DRAM[34523] = 8'b10001011;
DRAM[34524] = 8'b1111111;
DRAM[34525] = 8'b10010100;
DRAM[34526] = 8'b10010110;
DRAM[34527] = 8'b10010011;
DRAM[34528] = 8'b10001100;
DRAM[34529] = 8'b10010010;
DRAM[34530] = 8'b10001110;
DRAM[34531] = 8'b10000010;
DRAM[34532] = 8'b10000010;
DRAM[34533] = 8'b10001010;
DRAM[34534] = 8'b10000110;
DRAM[34535] = 8'b1111001;
DRAM[34536] = 8'b10000001;
DRAM[34537] = 8'b10000001;
DRAM[34538] = 8'b10000000;
DRAM[34539] = 8'b10000000;
DRAM[34540] = 8'b10000000;
DRAM[34541] = 8'b1111111;
DRAM[34542] = 8'b1111111;
DRAM[34543] = 8'b1111111;
DRAM[34544] = 8'b1111111;
DRAM[34545] = 8'b1111111;
DRAM[34546] = 8'b1111110;
DRAM[34547] = 8'b1111101;
DRAM[34548] = 8'b1111011;
DRAM[34549] = 8'b1111010;
DRAM[34550] = 8'b1111001;
DRAM[34551] = 8'b1111001;
DRAM[34552] = 8'b1111010;
DRAM[34553] = 8'b1111001;
DRAM[34554] = 8'b1111000;
DRAM[34555] = 8'b1110111;
DRAM[34556] = 8'b1110111;
DRAM[34557] = 8'b1110111;
DRAM[34558] = 8'b1110111;
DRAM[34559] = 8'b1111000;
DRAM[34560] = 8'b10001101;
DRAM[34561] = 8'b10001110;
DRAM[34562] = 8'b10001111;
DRAM[34563] = 8'b10010000;
DRAM[34564] = 8'b10010010;
DRAM[34565] = 8'b10010011;
DRAM[34566] = 8'b10010101;
DRAM[34567] = 8'b10010101;
DRAM[34568] = 8'b10010001;
DRAM[34569] = 8'b10010010;
DRAM[34570] = 8'b10010011;
DRAM[34571] = 8'b10010100;
DRAM[34572] = 8'b10010110;
DRAM[34573] = 8'b10010111;
DRAM[34574] = 8'b10011000;
DRAM[34575] = 8'b10011001;
DRAM[34576] = 8'b10011001;
DRAM[34577] = 8'b10011000;
DRAM[34578] = 8'b10011000;
DRAM[34579] = 8'b10011000;
DRAM[34580] = 8'b10011000;
DRAM[34581] = 8'b10011000;
DRAM[34582] = 8'b10011000;
DRAM[34583] = 8'b10011000;
DRAM[34584] = 8'b10011001;
DRAM[34585] = 8'b10011001;
DRAM[34586] = 8'b10011010;
DRAM[34587] = 8'b10011010;
DRAM[34588] = 8'b10011010;
DRAM[34589] = 8'b10011011;
DRAM[34590] = 8'b10011011;
DRAM[34591] = 8'b10011011;
DRAM[34592] = 8'b10011011;
DRAM[34593] = 8'b10011011;
DRAM[34594] = 8'b10011011;
DRAM[34595] = 8'b10011011;
DRAM[34596] = 8'b10011011;
DRAM[34597] = 8'b10011011;
DRAM[34598] = 8'b10011011;
DRAM[34599] = 8'b10011011;
DRAM[34600] = 8'b10011101;
DRAM[34601] = 8'b10011101;
DRAM[34602] = 8'b10011101;
DRAM[34603] = 8'b10011110;
DRAM[34604] = 8'b10011110;
DRAM[34605] = 8'b10011111;
DRAM[34606] = 8'b10100000;
DRAM[34607] = 8'b10100001;
DRAM[34608] = 8'b10011100;
DRAM[34609] = 8'b10101000;
DRAM[34610] = 8'b10100011;
DRAM[34611] = 8'b10100100;
DRAM[34612] = 8'b10100100;
DRAM[34613] = 8'b10101110;
DRAM[34614] = 8'b10111111;
DRAM[34615] = 8'b11000010;
DRAM[34616] = 8'b10111100;
DRAM[34617] = 8'b10110100;
DRAM[34618] = 8'b10110111;
DRAM[34619] = 8'b10101000;
DRAM[34620] = 8'b10101110;
DRAM[34621] = 8'b10001100;
DRAM[34622] = 8'b10010011;
DRAM[34623] = 8'b10100010;
DRAM[34624] = 8'b10111100;
DRAM[34625] = 8'b10111001;
DRAM[34626] = 8'b10101110;
DRAM[34627] = 8'b10100001;
DRAM[34628] = 8'b10011101;
DRAM[34629] = 8'b10011110;
DRAM[34630] = 8'b10011011;
DRAM[34631] = 8'b10010101;
DRAM[34632] = 8'b10001010;
DRAM[34633] = 8'b10001000;
DRAM[34634] = 8'b10000100;
DRAM[34635] = 8'b10000000;
DRAM[34636] = 8'b1111101;
DRAM[34637] = 8'b1111011;
DRAM[34638] = 8'b1111010;
DRAM[34639] = 8'b1111010;
DRAM[34640] = 8'b1111001;
DRAM[34641] = 8'b1111110;
DRAM[34642] = 8'b10001100;
DRAM[34643] = 8'b10011100;
DRAM[34644] = 8'b10100111;
DRAM[34645] = 8'b10101100;
DRAM[34646] = 8'b10110011;
DRAM[34647] = 8'b10111010;
DRAM[34648] = 8'b10110111;
DRAM[34649] = 8'b10101111;
DRAM[34650] = 8'b10101010;
DRAM[34651] = 8'b10101110;
DRAM[34652] = 8'b10110001;
DRAM[34653] = 8'b10101111;
DRAM[34654] = 8'b10101100;
DRAM[34655] = 8'b10101100;
DRAM[34656] = 8'b10100001;
DRAM[34657] = 8'b10100000;
DRAM[34658] = 8'b10100100;
DRAM[34659] = 8'b10101010;
DRAM[34660] = 8'b10101000;
DRAM[34661] = 8'b10100010;
DRAM[34662] = 8'b10100100;
DRAM[34663] = 8'b10101100;
DRAM[34664] = 8'b10000010;
DRAM[34665] = 8'b10100011;
DRAM[34666] = 8'b10011011;
DRAM[34667] = 8'b10110000;
DRAM[34668] = 8'b10010111;
DRAM[34669] = 8'b10010100;
DRAM[34670] = 8'b10100011;
DRAM[34671] = 8'b10101001;
DRAM[34672] = 8'b10011000;
DRAM[34673] = 8'b10100110;
DRAM[34674] = 8'b10111110;
DRAM[34675] = 8'b10111011;
DRAM[34676] = 8'b11001100;
DRAM[34677] = 8'b11001001;
DRAM[34678] = 8'b11001110;
DRAM[34679] = 8'b11000000;
DRAM[34680] = 8'b11000110;
DRAM[34681] = 8'b11011110;
DRAM[34682] = 8'b11101010;
DRAM[34683] = 8'b11100000;
DRAM[34684] = 8'b11011010;
DRAM[34685] = 8'b11100011;
DRAM[34686] = 8'b11101010;
DRAM[34687] = 8'b11101001;
DRAM[34688] = 8'b11111010;
DRAM[34689] = 8'b11111010;
DRAM[34690] = 8'b11111010;
DRAM[34691] = 8'b11111010;
DRAM[34692] = 8'b11111010;
DRAM[34693] = 8'b11111010;
DRAM[34694] = 8'b11111011;
DRAM[34695] = 8'b11111100;
DRAM[34696] = 8'b11111111;
DRAM[34697] = 8'b11111110;
DRAM[34698] = 8'b11111110;
DRAM[34699] = 8'b11111111;
DRAM[34700] = 8'b11111111;
DRAM[34701] = 8'b11111010;
DRAM[34702] = 8'b11111011;
DRAM[34703] = 8'b11111111;
DRAM[34704] = 8'b11111101;
DRAM[34705] = 8'b11111101;
DRAM[34706] = 8'b11111101;
DRAM[34707] = 8'b11111101;
DRAM[34708] = 8'b11111101;
DRAM[34709] = 8'b11111100;
DRAM[34710] = 8'b11111010;
DRAM[34711] = 8'b11111010;
DRAM[34712] = 8'b11111000;
DRAM[34713] = 8'b11110111;
DRAM[34714] = 8'b11110110;
DRAM[34715] = 8'b11111000;
DRAM[34716] = 8'b11111010;
DRAM[34717] = 8'b11111011;
DRAM[34718] = 8'b11111011;
DRAM[34719] = 8'b11111001;
DRAM[34720] = 8'b11111100;
DRAM[34721] = 8'b11111011;
DRAM[34722] = 8'b11111011;
DRAM[34723] = 8'b11111100;
DRAM[34724] = 8'b11111100;
DRAM[34725] = 8'b11111010;
DRAM[34726] = 8'b11110110;
DRAM[34727] = 8'b11110011;
DRAM[34728] = 8'b11111011;
DRAM[34729] = 8'b11011011;
DRAM[34730] = 8'b11010010;
DRAM[34731] = 8'b11011110;
DRAM[34732] = 8'b11011001;
DRAM[34733] = 8'b11001010;
DRAM[34734] = 8'b11000011;
DRAM[34735] = 8'b11000001;
DRAM[34736] = 8'b11010110;
DRAM[34737] = 8'b10110010;
DRAM[34738] = 8'b10101100;
DRAM[34739] = 8'b10110011;
DRAM[34740] = 8'b10100100;
DRAM[34741] = 8'b10011011;
DRAM[34742] = 8'b10100100;
DRAM[34743] = 8'b10100110;
DRAM[34744] = 8'b10101011;
DRAM[34745] = 8'b10101111;
DRAM[34746] = 8'b10101111;
DRAM[34747] = 8'b10101100;
DRAM[34748] = 8'b10101101;
DRAM[34749] = 8'b10101111;
DRAM[34750] = 8'b10101010;
DRAM[34751] = 8'b10100001;
DRAM[34752] = 8'b10011101;
DRAM[34753] = 8'b10010001;
DRAM[34754] = 8'b10000101;
DRAM[34755] = 8'b10000011;
DRAM[34756] = 8'b10000111;
DRAM[34757] = 8'b10001100;
DRAM[34758] = 8'b10010010;
DRAM[34759] = 8'b10011000;
DRAM[34760] = 8'b10100100;
DRAM[34761] = 8'b10110011;
DRAM[34762] = 8'b11001001;
DRAM[34763] = 8'b11100001;
DRAM[34764] = 8'b11110010;
DRAM[34765] = 8'b11110011;
DRAM[34766] = 8'b11100001;
DRAM[34767] = 8'b11001101;
DRAM[34768] = 8'b10110100;
DRAM[34769] = 8'b10010010;
DRAM[34770] = 8'b10000110;
DRAM[34771] = 8'b10010010;
DRAM[34772] = 8'b10001111;
DRAM[34773] = 8'b10000111;
DRAM[34774] = 8'b10001101;
DRAM[34775] = 8'b10010110;
DRAM[34776] = 8'b10000000;
DRAM[34777] = 8'b10011010;
DRAM[34778] = 8'b10010000;
DRAM[34779] = 8'b10011001;
DRAM[34780] = 8'b1110101;
DRAM[34781] = 8'b10011001;
DRAM[34782] = 8'b10000101;
DRAM[34783] = 8'b1110101;
DRAM[34784] = 8'b10000111;
DRAM[34785] = 8'b10100001;
DRAM[34786] = 8'b10101000;
DRAM[34787] = 8'b10001111;
DRAM[34788] = 8'b1111100;
DRAM[34789] = 8'b10000000;
DRAM[34790] = 8'b10000110;
DRAM[34791] = 8'b10000100;
DRAM[34792] = 8'b10000001;
DRAM[34793] = 8'b10000001;
DRAM[34794] = 8'b10000001;
DRAM[34795] = 8'b10000000;
DRAM[34796] = 8'b10000000;
DRAM[34797] = 8'b1111111;
DRAM[34798] = 8'b1111111;
DRAM[34799] = 8'b1111111;
DRAM[34800] = 8'b10000000;
DRAM[34801] = 8'b1111111;
DRAM[34802] = 8'b1111110;
DRAM[34803] = 8'b1111101;
DRAM[34804] = 8'b1111011;
DRAM[34805] = 8'b1111010;
DRAM[34806] = 8'b1111001;
DRAM[34807] = 8'b1111001;
DRAM[34808] = 8'b1111010;
DRAM[34809] = 8'b1111001;
DRAM[34810] = 8'b1111000;
DRAM[34811] = 8'b1110111;
DRAM[34812] = 8'b1110111;
DRAM[34813] = 8'b1110111;
DRAM[34814] = 8'b1110111;
DRAM[34815] = 8'b1111000;
DRAM[34816] = 8'b10001101;
DRAM[34817] = 8'b10001111;
DRAM[34818] = 8'b10010010;
DRAM[34819] = 8'b10010101;
DRAM[34820] = 8'b10010110;
DRAM[34821] = 8'b10010110;
DRAM[34822] = 8'b10010101;
DRAM[34823] = 8'b10010100;
DRAM[34824] = 8'b10010011;
DRAM[34825] = 8'b10010100;
DRAM[34826] = 8'b10010100;
DRAM[34827] = 8'b10010101;
DRAM[34828] = 8'b10010110;
DRAM[34829] = 8'b10010111;
DRAM[34830] = 8'b10011000;
DRAM[34831] = 8'b10011000;
DRAM[34832] = 8'b10010101;
DRAM[34833] = 8'b10010110;
DRAM[34834] = 8'b10010111;
DRAM[34835] = 8'b10011000;
DRAM[34836] = 8'b10011001;
DRAM[34837] = 8'b10011001;
DRAM[34838] = 8'b10011001;
DRAM[34839] = 8'b10011001;
DRAM[34840] = 8'b10011000;
DRAM[34841] = 8'b10011000;
DRAM[34842] = 8'b10011001;
DRAM[34843] = 8'b10011001;
DRAM[34844] = 8'b10011010;
DRAM[34845] = 8'b10011011;
DRAM[34846] = 8'b10011100;
DRAM[34847] = 8'b10011100;
DRAM[34848] = 8'b10011010;
DRAM[34849] = 8'b10011011;
DRAM[34850] = 8'b10011011;
DRAM[34851] = 8'b10011100;
DRAM[34852] = 8'b10011101;
DRAM[34853] = 8'b10011110;
DRAM[34854] = 8'b10011111;
DRAM[34855] = 8'b10011111;
DRAM[34856] = 8'b10011110;
DRAM[34857] = 8'b10011110;
DRAM[34858] = 8'b10011110;
DRAM[34859] = 8'b10011110;
DRAM[34860] = 8'b10011110;
DRAM[34861] = 8'b10011110;
DRAM[34862] = 8'b10011110;
DRAM[34863] = 8'b10011110;
DRAM[34864] = 8'b10011001;
DRAM[34865] = 8'b10011001;
DRAM[34866] = 8'b10011110;
DRAM[34867] = 8'b10100101;
DRAM[34868] = 8'b10101011;
DRAM[34869] = 8'b10110011;
DRAM[34870] = 8'b11000000;
DRAM[34871] = 8'b11001101;
DRAM[34872] = 8'b11001101;
DRAM[34873] = 8'b10111100;
DRAM[34874] = 8'b10110110;
DRAM[34875] = 8'b10110101;
DRAM[34876] = 8'b10011110;
DRAM[34877] = 8'b10000110;
DRAM[34878] = 8'b10010111;
DRAM[34879] = 8'b10111111;
DRAM[34880] = 8'b11000110;
DRAM[34881] = 8'b10111010;
DRAM[34882] = 8'b10101110;
DRAM[34883] = 8'b10101001;
DRAM[34884] = 8'b10100110;
DRAM[34885] = 8'b10100001;
DRAM[34886] = 8'b10011111;
DRAM[34887] = 8'b10100000;
DRAM[34888] = 8'b10011100;
DRAM[34889] = 8'b10010101;
DRAM[34890] = 8'b10001100;
DRAM[34891] = 8'b10001001;
DRAM[34892] = 8'b10001001;
DRAM[34893] = 8'b10001000;
DRAM[34894] = 8'b10000010;
DRAM[34895] = 8'b1111101;
DRAM[34896] = 8'b1111100;
DRAM[34897] = 8'b1111110;
DRAM[34898] = 8'b10000111;
DRAM[34899] = 8'b10010101;
DRAM[34900] = 8'b10100010;
DRAM[34901] = 8'b10100111;
DRAM[34902] = 8'b10100110;
DRAM[34903] = 8'b10100101;
DRAM[34904] = 8'b10101101;
DRAM[34905] = 8'b10101111;
DRAM[34906] = 8'b10110011;
DRAM[34907] = 8'b10110110;
DRAM[34908] = 8'b10110101;
DRAM[34909] = 8'b10110010;
DRAM[34910] = 8'b10101100;
DRAM[34911] = 8'b10101000;
DRAM[34912] = 8'b10101010;
DRAM[34913] = 8'b10011001;
DRAM[34914] = 8'b10010100;
DRAM[34915] = 8'b10100000;
DRAM[34916] = 8'b10100111;
DRAM[34917] = 8'b10011111;
DRAM[34918] = 8'b10011001;
DRAM[34919] = 8'b10011011;
DRAM[34920] = 8'b10100111;
DRAM[34921] = 8'b10100111;
DRAM[34922] = 8'b10110110;
DRAM[34923] = 8'b10011100;
DRAM[34924] = 8'b1110111;
DRAM[34925] = 8'b10011010;
DRAM[34926] = 8'b10111000;
DRAM[34927] = 8'b10010001;
DRAM[34928] = 8'b10101111;
DRAM[34929] = 8'b10110000;
DRAM[34930] = 8'b10111001;
DRAM[34931] = 8'b11000111;
DRAM[34932] = 8'b11001001;
DRAM[34933] = 8'b11000001;
DRAM[34934] = 8'b10111110;
DRAM[34935] = 8'b11000010;
DRAM[34936] = 8'b11011100;
DRAM[34937] = 8'b11011100;
DRAM[34938] = 8'b11011110;
DRAM[34939] = 8'b11100001;
DRAM[34940] = 8'b11100111;
DRAM[34941] = 8'b11101111;
DRAM[34942] = 8'b11110110;
DRAM[34943] = 8'b11111010;
DRAM[34944] = 8'b11110110;
DRAM[34945] = 8'b11111011;
DRAM[34946] = 8'b11111101;
DRAM[34947] = 8'b11111010;
DRAM[34948] = 8'b11111010;
DRAM[34949] = 8'b11111110;
DRAM[34950] = 8'b11111101;
DRAM[34951] = 8'b11110111;
DRAM[34952] = 8'b11111101;
DRAM[34953] = 8'b11111101;
DRAM[34954] = 8'b11111110;
DRAM[34955] = 8'b11111110;
DRAM[34956] = 8'b11111110;
DRAM[34957] = 8'b11111101;
DRAM[34958] = 8'b11111100;
DRAM[34959] = 8'b11111100;
DRAM[34960] = 8'b11111101;
DRAM[34961] = 8'b11111101;
DRAM[34962] = 8'b11111101;
DRAM[34963] = 8'b11111111;
DRAM[34964] = 8'b11111111;
DRAM[34965] = 8'b11111111;
DRAM[34966] = 8'b11111101;
DRAM[34967] = 8'b11111011;
DRAM[34968] = 8'b11111010;
DRAM[34969] = 8'b11111001;
DRAM[34970] = 8'b11111001;
DRAM[34971] = 8'b11111000;
DRAM[34972] = 8'b11110111;
DRAM[34973] = 8'b11110111;
DRAM[34974] = 8'b11110110;
DRAM[34975] = 8'b11110110;
DRAM[34976] = 8'b11110011;
DRAM[34977] = 8'b11111000;
DRAM[34978] = 8'b11111100;
DRAM[34979] = 8'b11111100;
DRAM[34980] = 8'b11111010;
DRAM[34981] = 8'b11110111;
DRAM[34982] = 8'b11110011;
DRAM[34983] = 8'b11110000;
DRAM[34984] = 8'b11101100;
DRAM[34985] = 8'b11101110;
DRAM[34986] = 8'b11100010;
DRAM[34987] = 8'b11010000;
DRAM[34988] = 8'b11010011;
DRAM[34989] = 8'b11011101;
DRAM[34990] = 8'b11010001;
DRAM[34991] = 8'b10110111;
DRAM[34992] = 8'b10110010;
DRAM[34993] = 8'b10110111;
DRAM[34994] = 8'b10111010;
DRAM[34995] = 8'b10111000;
DRAM[34996] = 8'b10110001;
DRAM[34997] = 8'b10110000;
DRAM[34998] = 8'b10110110;
DRAM[34999] = 8'b10111110;
DRAM[35000] = 8'b10111010;
DRAM[35001] = 8'b10111000;
DRAM[35002] = 8'b10111000;
DRAM[35003] = 8'b10111000;
DRAM[35004] = 8'b10111000;
DRAM[35005] = 8'b10110100;
DRAM[35006] = 8'b10101011;
DRAM[35007] = 8'b10100100;
DRAM[35008] = 8'b10010000;
DRAM[35009] = 8'b10001010;
DRAM[35010] = 8'b10000100;
DRAM[35011] = 8'b10000010;
DRAM[35012] = 8'b10000001;
DRAM[35013] = 8'b10000110;
DRAM[35014] = 8'b10010100;
DRAM[35015] = 8'b10100001;
DRAM[35016] = 8'b10101000;
DRAM[35017] = 8'b10110110;
DRAM[35018] = 8'b11001100;
DRAM[35019] = 8'b11100011;
DRAM[35020] = 8'b11110100;
DRAM[35021] = 8'b11110100;
DRAM[35022] = 8'b11100000;
DRAM[35023] = 8'b11001011;
DRAM[35024] = 8'b10110011;
DRAM[35025] = 8'b10011101;
DRAM[35026] = 8'b10001101;
DRAM[35027] = 8'b10001110;
DRAM[35028] = 8'b10001111;
DRAM[35029] = 8'b10000111;
DRAM[35030] = 8'b10000101;
DRAM[35031] = 8'b10001100;
DRAM[35032] = 8'b10001001;
DRAM[35033] = 8'b10001001;
DRAM[35034] = 8'b10001000;
DRAM[35035] = 8'b10001000;
DRAM[35036] = 8'b10001000;
DRAM[35037] = 8'b10001001;
DRAM[35038] = 8'b10001010;
DRAM[35039] = 8'b10001010;
DRAM[35040] = 8'b10000010;
DRAM[35041] = 8'b10000100;
DRAM[35042] = 8'b10000111;
DRAM[35043] = 8'b10001010;
DRAM[35044] = 8'b10001011;
DRAM[35045] = 8'b10001001;
DRAM[35046] = 8'b10000111;
DRAM[35047] = 8'b10000101;
DRAM[35048] = 8'b10000010;
DRAM[35049] = 8'b10000000;
DRAM[35050] = 8'b1111111;
DRAM[35051] = 8'b1111101;
DRAM[35052] = 8'b1111101;
DRAM[35053] = 8'b1111110;
DRAM[35054] = 8'b1111111;
DRAM[35055] = 8'b1111111;
DRAM[35056] = 8'b10000000;
DRAM[35057] = 8'b1111111;
DRAM[35058] = 8'b1111110;
DRAM[35059] = 8'b1111101;
DRAM[35060] = 8'b1111100;
DRAM[35061] = 8'b1111011;
DRAM[35062] = 8'b1111100;
DRAM[35063] = 8'b1111100;
DRAM[35064] = 8'b1111000;
DRAM[35065] = 8'b1111000;
DRAM[35066] = 8'b1111000;
DRAM[35067] = 8'b1110111;
DRAM[35068] = 8'b1110111;
DRAM[35069] = 8'b1110110;
DRAM[35070] = 8'b1110110;
DRAM[35071] = 8'b1110110;
DRAM[35072] = 8'b10001110;
DRAM[35073] = 8'b10010000;
DRAM[35074] = 8'b10010010;
DRAM[35075] = 8'b10010101;
DRAM[35076] = 8'b10010110;
DRAM[35077] = 8'b10010110;
DRAM[35078] = 8'b10010101;
DRAM[35079] = 8'b10010100;
DRAM[35080] = 8'b10010101;
DRAM[35081] = 8'b10010101;
DRAM[35082] = 8'b10010110;
DRAM[35083] = 8'b10010110;
DRAM[35084] = 8'b10010111;
DRAM[35085] = 8'b10011000;
DRAM[35086] = 8'b10011001;
DRAM[35087] = 8'b10011001;
DRAM[35088] = 8'b10011001;
DRAM[35089] = 8'b10011001;
DRAM[35090] = 8'b10011010;
DRAM[35091] = 8'b10011011;
DRAM[35092] = 8'b10011011;
DRAM[35093] = 8'b10011011;
DRAM[35094] = 8'b10011010;
DRAM[35095] = 8'b10011010;
DRAM[35096] = 8'b10011000;
DRAM[35097] = 8'b10011001;
DRAM[35098] = 8'b10011001;
DRAM[35099] = 8'b10011010;
DRAM[35100] = 8'b10011011;
DRAM[35101] = 8'b10011100;
DRAM[35102] = 8'b10011100;
DRAM[35103] = 8'b10011100;
DRAM[35104] = 8'b10011100;
DRAM[35105] = 8'b10011100;
DRAM[35106] = 8'b10011101;
DRAM[35107] = 8'b10011101;
DRAM[35108] = 8'b10011110;
DRAM[35109] = 8'b10011110;
DRAM[35110] = 8'b10011111;
DRAM[35111] = 8'b10011111;
DRAM[35112] = 8'b10011111;
DRAM[35113] = 8'b10011111;
DRAM[35114] = 8'b10011111;
DRAM[35115] = 8'b10011111;
DRAM[35116] = 8'b10011111;
DRAM[35117] = 8'b10011111;
DRAM[35118] = 8'b10011111;
DRAM[35119] = 8'b10011111;
DRAM[35120] = 8'b10100110;
DRAM[35121] = 8'b10100100;
DRAM[35122] = 8'b10100011;
DRAM[35123] = 8'b10100101;
DRAM[35124] = 8'b10100110;
DRAM[35125] = 8'b10101010;
DRAM[35126] = 8'b10110100;
DRAM[35127] = 8'b11000000;
DRAM[35128] = 8'b11010101;
DRAM[35129] = 8'b10111101;
DRAM[35130] = 8'b10101100;
DRAM[35131] = 8'b10101010;
DRAM[35132] = 8'b10100100;
DRAM[35133] = 8'b10100011;
DRAM[35134] = 8'b10111011;
DRAM[35135] = 8'b11011101;
DRAM[35136] = 8'b11001000;
DRAM[35137] = 8'b10111101;
DRAM[35138] = 8'b10110001;
DRAM[35139] = 8'b10101011;
DRAM[35140] = 8'b10100111;
DRAM[35141] = 8'b10100001;
DRAM[35142] = 8'b10011101;
DRAM[35143] = 8'b10011101;
DRAM[35144] = 8'b10010111;
DRAM[35145] = 8'b10010100;
DRAM[35146] = 8'b10001111;
DRAM[35147] = 8'b10001001;
DRAM[35148] = 8'b10000101;
DRAM[35149] = 8'b10000010;
DRAM[35150] = 8'b10000000;
DRAM[35151] = 8'b1111110;
DRAM[35152] = 8'b1110101;
DRAM[35153] = 8'b1111110;
DRAM[35154] = 8'b10001010;
DRAM[35155] = 8'b10010101;
DRAM[35156] = 8'b10011010;
DRAM[35157] = 8'b10011100;
DRAM[35158] = 8'b10011110;
DRAM[35159] = 8'b10100001;
DRAM[35160] = 8'b10101110;
DRAM[35161] = 8'b10110001;
DRAM[35162] = 8'b10110100;
DRAM[35163] = 8'b10110110;
DRAM[35164] = 8'b10110101;
DRAM[35165] = 8'b10110011;
DRAM[35166] = 8'b10110010;
DRAM[35167] = 8'b10110010;
DRAM[35168] = 8'b10110010;
DRAM[35169] = 8'b10101001;
DRAM[35170] = 8'b10100101;
DRAM[35171] = 8'b10101010;
DRAM[35172] = 8'b10101011;
DRAM[35173] = 8'b10100101;
DRAM[35174] = 8'b10100011;
DRAM[35175] = 8'b10100101;
DRAM[35176] = 8'b10100110;
DRAM[35177] = 8'b10101100;
DRAM[35178] = 8'b10110000;
DRAM[35179] = 8'b10100010;
DRAM[35180] = 8'b10010100;
DRAM[35181] = 8'b10011101;
DRAM[35182] = 8'b10100100;
DRAM[35183] = 8'b10010110;
DRAM[35184] = 8'b10101100;
DRAM[35185] = 8'b10111010;
DRAM[35186] = 8'b11000111;
DRAM[35187] = 8'b11001001;
DRAM[35188] = 8'b11000111;
DRAM[35189] = 8'b11000111;
DRAM[35190] = 8'b11001001;
DRAM[35191] = 8'b11001010;
DRAM[35192] = 8'b11010111;
DRAM[35193] = 8'b11011100;
DRAM[35194] = 8'b11100011;
DRAM[35195] = 8'b11101010;
DRAM[35196] = 8'b11110000;
DRAM[35197] = 8'b11110011;
DRAM[35198] = 8'b11110100;
DRAM[35199] = 8'b11110100;
DRAM[35200] = 8'b11110101;
DRAM[35201] = 8'b11111001;
DRAM[35202] = 8'b11111010;
DRAM[35203] = 8'b11110110;
DRAM[35204] = 8'b11110110;
DRAM[35205] = 8'b11111001;
DRAM[35206] = 8'b11111001;
DRAM[35207] = 8'b11110100;
DRAM[35208] = 8'b11111101;
DRAM[35209] = 8'b11111101;
DRAM[35210] = 8'b11111110;
DRAM[35211] = 8'b11111101;
DRAM[35212] = 8'b11111101;
DRAM[35213] = 8'b11111100;
DRAM[35214] = 8'b11111011;
DRAM[35215] = 8'b11111010;
DRAM[35216] = 8'b11111011;
DRAM[35217] = 8'b11111010;
DRAM[35218] = 8'b11111001;
DRAM[35219] = 8'b11111010;
DRAM[35220] = 8'b11111011;
DRAM[35221] = 8'b11111100;
DRAM[35222] = 8'b11111010;
DRAM[35223] = 8'b11111000;
DRAM[35224] = 8'b11110110;
DRAM[35225] = 8'b11110101;
DRAM[35226] = 8'b11110011;
DRAM[35227] = 8'b11110001;
DRAM[35228] = 8'b11110001;
DRAM[35229] = 8'b11110010;
DRAM[35230] = 8'b11110100;
DRAM[35231] = 8'b11110110;
DRAM[35232] = 8'b11110110;
DRAM[35233] = 8'b11111000;
DRAM[35234] = 8'b11111001;
DRAM[35235] = 8'b11110111;
DRAM[35236] = 8'b11110101;
DRAM[35237] = 8'b11110100;
DRAM[35238] = 8'b11110011;
DRAM[35239] = 8'b11110010;
DRAM[35240] = 8'b11110100;
DRAM[35241] = 8'b11110101;
DRAM[35242] = 8'b11101010;
DRAM[35243] = 8'b11011010;
DRAM[35244] = 8'b11010111;
DRAM[35245] = 8'b11011101;
DRAM[35246] = 8'b11010110;
DRAM[35247] = 8'b11000110;
DRAM[35248] = 8'b10111111;
DRAM[35249] = 8'b11000010;
DRAM[35250] = 8'b10111000;
DRAM[35251] = 8'b10100111;
DRAM[35252] = 8'b10101001;
DRAM[35253] = 8'b10111001;
DRAM[35254] = 8'b10111010;
DRAM[35255] = 8'b10101101;
DRAM[35256] = 8'b11000100;
DRAM[35257] = 8'b10111110;
DRAM[35258] = 8'b10110110;
DRAM[35259] = 8'b10101111;
DRAM[35260] = 8'b10101010;
DRAM[35261] = 8'b10100010;
DRAM[35262] = 8'b10011001;
DRAM[35263] = 8'b10010011;
DRAM[35264] = 8'b10000111;
DRAM[35265] = 8'b10000101;
DRAM[35266] = 8'b10000110;
DRAM[35267] = 8'b10001010;
DRAM[35268] = 8'b10001101;
DRAM[35269] = 8'b10001110;
DRAM[35270] = 8'b10010011;
DRAM[35271] = 8'b10011010;
DRAM[35272] = 8'b10101011;
DRAM[35273] = 8'b11000000;
DRAM[35274] = 8'b11011011;
DRAM[35275] = 8'b11101111;
DRAM[35276] = 8'b11110111;
DRAM[35277] = 8'b11110010;
DRAM[35278] = 8'b11100010;
DRAM[35279] = 8'b11010011;
DRAM[35280] = 8'b10101010;
DRAM[35281] = 8'b10011011;
DRAM[35282] = 8'b10010001;
DRAM[35283] = 8'b10010001;
DRAM[35284] = 8'b10010001;
DRAM[35285] = 8'b10001100;
DRAM[35286] = 8'b10001010;
DRAM[35287] = 8'b10001101;
DRAM[35288] = 8'b10001010;
DRAM[35289] = 8'b10001001;
DRAM[35290] = 8'b10001001;
DRAM[35291] = 8'b10001000;
DRAM[35292] = 8'b10001000;
DRAM[35293] = 8'b10001001;
DRAM[35294] = 8'b10001010;
DRAM[35295] = 8'b10001010;
DRAM[35296] = 8'b10000101;
DRAM[35297] = 8'b10000110;
DRAM[35298] = 8'b10001000;
DRAM[35299] = 8'b10001000;
DRAM[35300] = 8'b10000111;
DRAM[35301] = 8'b10000110;
DRAM[35302] = 8'b10000011;
DRAM[35303] = 8'b10000010;
DRAM[35304] = 8'b10000001;
DRAM[35305] = 8'b10000001;
DRAM[35306] = 8'b10000000;
DRAM[35307] = 8'b1111111;
DRAM[35308] = 8'b1111111;
DRAM[35309] = 8'b1111111;
DRAM[35310] = 8'b1111111;
DRAM[35311] = 8'b1111111;
DRAM[35312] = 8'b10000000;
DRAM[35313] = 8'b1111111;
DRAM[35314] = 8'b1111110;
DRAM[35315] = 8'b1111101;
DRAM[35316] = 8'b1111100;
DRAM[35317] = 8'b1111011;
DRAM[35318] = 8'b1111100;
DRAM[35319] = 8'b1111100;
DRAM[35320] = 8'b1111000;
DRAM[35321] = 8'b1111000;
DRAM[35322] = 8'b1111000;
DRAM[35323] = 8'b1110111;
DRAM[35324] = 8'b1110111;
DRAM[35325] = 8'b1110111;
DRAM[35326] = 8'b1110110;
DRAM[35327] = 8'b1110110;
DRAM[35328] = 8'b10001111;
DRAM[35329] = 8'b10010001;
DRAM[35330] = 8'b10010011;
DRAM[35331] = 8'b10010101;
DRAM[35332] = 8'b10010111;
DRAM[35333] = 8'b10010111;
DRAM[35334] = 8'b10010110;
DRAM[35335] = 8'b10010110;
DRAM[35336] = 8'b10010111;
DRAM[35337] = 8'b10010111;
DRAM[35338] = 8'b10011000;
DRAM[35339] = 8'b10011000;
DRAM[35340] = 8'b10011001;
DRAM[35341] = 8'b10011010;
DRAM[35342] = 8'b10011010;
DRAM[35343] = 8'b10011011;
DRAM[35344] = 8'b10011100;
DRAM[35345] = 8'b10011101;
DRAM[35346] = 8'b10011101;
DRAM[35347] = 8'b10011101;
DRAM[35348] = 8'b10011101;
DRAM[35349] = 8'b10011100;
DRAM[35350] = 8'b10011100;
DRAM[35351] = 8'b10011011;
DRAM[35352] = 8'b10011001;
DRAM[35353] = 8'b10011001;
DRAM[35354] = 8'b10011010;
DRAM[35355] = 8'b10011011;
DRAM[35356] = 8'b10011100;
DRAM[35357] = 8'b10011100;
DRAM[35358] = 8'b10011101;
DRAM[35359] = 8'b10011101;
DRAM[35360] = 8'b10011110;
DRAM[35361] = 8'b10011110;
DRAM[35362] = 8'b10011110;
DRAM[35363] = 8'b10011111;
DRAM[35364] = 8'b10011111;
DRAM[35365] = 8'b10011111;
DRAM[35366] = 8'b10011111;
DRAM[35367] = 8'b10011111;
DRAM[35368] = 8'b10100001;
DRAM[35369] = 8'b10100001;
DRAM[35370] = 8'b10100001;
DRAM[35371] = 8'b10100001;
DRAM[35372] = 8'b10100001;
DRAM[35373] = 8'b10100001;
DRAM[35374] = 8'b10100001;
DRAM[35375] = 8'b10100001;
DRAM[35376] = 8'b10100100;
DRAM[35377] = 8'b10100001;
DRAM[35378] = 8'b10100000;
DRAM[35379] = 8'b10100001;
DRAM[35380] = 8'b10100010;
DRAM[35381] = 8'b10100111;
DRAM[35382] = 8'b10110011;
DRAM[35383] = 8'b11000000;
DRAM[35384] = 8'b11000111;
DRAM[35385] = 8'b10111010;
DRAM[35386] = 8'b10110011;
DRAM[35387] = 8'b10111100;
DRAM[35388] = 8'b11001001;
DRAM[35389] = 8'b11010010;
DRAM[35390] = 8'b11011010;
DRAM[35391] = 8'b11100001;
DRAM[35392] = 8'b11001011;
DRAM[35393] = 8'b10111111;
DRAM[35394] = 8'b10110100;
DRAM[35395] = 8'b10101111;
DRAM[35396] = 8'b10101010;
DRAM[35397] = 8'b10100010;
DRAM[35398] = 8'b10011101;
DRAM[35399] = 8'b10011100;
DRAM[35400] = 8'b10011001;
DRAM[35401] = 8'b10011001;
DRAM[35402] = 8'b10010101;
DRAM[35403] = 8'b10001111;
DRAM[35404] = 8'b10000111;
DRAM[35405] = 8'b10000011;
DRAM[35406] = 8'b10000010;
DRAM[35407] = 8'b10000011;
DRAM[35408] = 8'b1111100;
DRAM[35409] = 8'b10001010;
DRAM[35410] = 8'b10011010;
DRAM[35411] = 8'b10100000;
DRAM[35412] = 8'b10011101;
DRAM[35413] = 8'b10011100;
DRAM[35414] = 8'b10100001;
DRAM[35415] = 8'b10100111;
DRAM[35416] = 8'b10100100;
DRAM[35417] = 8'b10101010;
DRAM[35418] = 8'b10110010;
DRAM[35419] = 8'b10110101;
DRAM[35420] = 8'b10110100;
DRAM[35421] = 8'b10110001;
DRAM[35422] = 8'b10110000;
DRAM[35423] = 8'b10110000;
DRAM[35424] = 8'b10111110;
DRAM[35425] = 8'b10111010;
DRAM[35426] = 8'b10110011;
DRAM[35427] = 8'b10101010;
DRAM[35428] = 8'b10100001;
DRAM[35429] = 8'b10011001;
DRAM[35430] = 8'b10010101;
DRAM[35431] = 8'b10010100;
DRAM[35432] = 8'b10001110;
DRAM[35433] = 8'b10011000;
DRAM[35434] = 8'b10010011;
DRAM[35435] = 8'b10010100;
DRAM[35436] = 8'b10100010;
DRAM[35437] = 8'b10011101;
DRAM[35438] = 8'b10011010;
DRAM[35439] = 8'b10101011;
DRAM[35440] = 8'b10101100;
DRAM[35441] = 8'b11000010;
DRAM[35442] = 8'b11001111;
DRAM[35443] = 8'b11000111;
DRAM[35444] = 8'b10111111;
DRAM[35445] = 8'b11000100;
DRAM[35446] = 8'b11001100;
DRAM[35447] = 8'b11001101;
DRAM[35448] = 8'b11011010;
DRAM[35449] = 8'b11011111;
DRAM[35450] = 8'b11100110;
DRAM[35451] = 8'b11101110;
DRAM[35452] = 8'b11110011;
DRAM[35453] = 8'b11110100;
DRAM[35454] = 8'b11110100;
DRAM[35455] = 8'b11110011;
DRAM[35456] = 8'b11111010;
DRAM[35457] = 8'b11111100;
DRAM[35458] = 8'b11111010;
DRAM[35459] = 8'b11110111;
DRAM[35460] = 8'b11110110;
DRAM[35461] = 8'b11111000;
DRAM[35462] = 8'b11111000;
DRAM[35463] = 8'b11110110;
DRAM[35464] = 8'b11111010;
DRAM[35465] = 8'b11111010;
DRAM[35466] = 8'b11111010;
DRAM[35467] = 8'b11111010;
DRAM[35468] = 8'b11111010;
DRAM[35469] = 8'b11111001;
DRAM[35470] = 8'b11111000;
DRAM[35471] = 8'b11110111;
DRAM[35472] = 8'b11111010;
DRAM[35473] = 8'b11111001;
DRAM[35474] = 8'b11110111;
DRAM[35475] = 8'b11111000;
DRAM[35476] = 8'b11111010;
DRAM[35477] = 8'b11111010;
DRAM[35478] = 8'b11111001;
DRAM[35479] = 8'b11111000;
DRAM[35480] = 8'b11110110;
DRAM[35481] = 8'b11110101;
DRAM[35482] = 8'b11110010;
DRAM[35483] = 8'b11110000;
DRAM[35484] = 8'b11110001;
DRAM[35485] = 8'b11110011;
DRAM[35486] = 8'b11110110;
DRAM[35487] = 8'b11111000;
DRAM[35488] = 8'b11111011;
DRAM[35489] = 8'b11111001;
DRAM[35490] = 8'b11110111;
DRAM[35491] = 8'b11110110;
DRAM[35492] = 8'b11110110;
DRAM[35493] = 8'b11110111;
DRAM[35494] = 8'b11111001;
DRAM[35495] = 8'b11111011;
DRAM[35496] = 8'b11110011;
DRAM[35497] = 8'b11110011;
DRAM[35498] = 8'b11101100;
DRAM[35499] = 8'b11011111;
DRAM[35500] = 8'b11010101;
DRAM[35501] = 8'b11010001;
DRAM[35502] = 8'b11010000;
DRAM[35503] = 8'b11001110;
DRAM[35504] = 8'b11000100;
DRAM[35505] = 8'b10111000;
DRAM[35506] = 8'b10110110;
DRAM[35507] = 8'b10111111;
DRAM[35508] = 8'b10111011;
DRAM[35509] = 8'b10101110;
DRAM[35510] = 8'b10101110;
DRAM[35511] = 8'b10111011;
DRAM[35512] = 8'b10100100;
DRAM[35513] = 8'b10101011;
DRAM[35514] = 8'b10110111;
DRAM[35515] = 8'b11000010;
DRAM[35516] = 8'b11000100;
DRAM[35517] = 8'b10111010;
DRAM[35518] = 8'b10101000;
DRAM[35519] = 8'b10011001;
DRAM[35520] = 8'b10010101;
DRAM[35521] = 8'b10001100;
DRAM[35522] = 8'b10000100;
DRAM[35523] = 8'b10000100;
DRAM[35524] = 8'b10001000;
DRAM[35525] = 8'b10001111;
DRAM[35526] = 8'b10011001;
DRAM[35527] = 8'b10100010;
DRAM[35528] = 8'b10101011;
DRAM[35529] = 8'b10111110;
DRAM[35530] = 8'b11010101;
DRAM[35531] = 8'b11100101;
DRAM[35532] = 8'b11101001;
DRAM[35533] = 8'b11100000;
DRAM[35534] = 8'b11001010;
DRAM[35535] = 8'b10110111;
DRAM[35536] = 8'b10011010;
DRAM[35537] = 8'b10010110;
DRAM[35538] = 8'b10010010;
DRAM[35539] = 8'b10010001;
DRAM[35540] = 8'b10010000;
DRAM[35541] = 8'b10010000;
DRAM[35542] = 8'b10001110;
DRAM[35543] = 8'b10001100;
DRAM[35544] = 8'b10001011;
DRAM[35545] = 8'b10001010;
DRAM[35546] = 8'b10001010;
DRAM[35547] = 8'b10001001;
DRAM[35548] = 8'b10001001;
DRAM[35549] = 8'b10001001;
DRAM[35550] = 8'b10001010;
DRAM[35551] = 8'b10001010;
DRAM[35552] = 8'b10001010;
DRAM[35553] = 8'b10001001;
DRAM[35554] = 8'b10001000;
DRAM[35555] = 8'b10000110;
DRAM[35556] = 8'b10000100;
DRAM[35557] = 8'b10000010;
DRAM[35558] = 8'b10000000;
DRAM[35559] = 8'b1111111;
DRAM[35560] = 8'b10000001;
DRAM[35561] = 8'b10000001;
DRAM[35562] = 8'b10000010;
DRAM[35563] = 8'b10000010;
DRAM[35564] = 8'b10000001;
DRAM[35565] = 8'b10000001;
DRAM[35566] = 8'b10000000;
DRAM[35567] = 8'b1111111;
DRAM[35568] = 8'b10000000;
DRAM[35569] = 8'b1111111;
DRAM[35570] = 8'b1111110;
DRAM[35571] = 8'b1111101;
DRAM[35572] = 8'b1111100;
DRAM[35573] = 8'b1111011;
DRAM[35574] = 8'b1111100;
DRAM[35575] = 8'b1111100;
DRAM[35576] = 8'b1111000;
DRAM[35577] = 8'b1111000;
DRAM[35578] = 8'b1111000;
DRAM[35579] = 8'b1111000;
DRAM[35580] = 8'b1110111;
DRAM[35581] = 8'b1110111;
DRAM[35582] = 8'b1110111;
DRAM[35583] = 8'b1110110;
DRAM[35584] = 8'b10010001;
DRAM[35585] = 8'b10010010;
DRAM[35586] = 8'b10010100;
DRAM[35587] = 8'b10010110;
DRAM[35588] = 8'b10010111;
DRAM[35589] = 8'b10011000;
DRAM[35590] = 8'b10011000;
DRAM[35591] = 8'b10010111;
DRAM[35592] = 8'b10011001;
DRAM[35593] = 8'b10011001;
DRAM[35594] = 8'b10011010;
DRAM[35595] = 8'b10011010;
DRAM[35596] = 8'b10011011;
DRAM[35597] = 8'b10011011;
DRAM[35598] = 8'b10011100;
DRAM[35599] = 8'b10011100;
DRAM[35600] = 8'b10011110;
DRAM[35601] = 8'b10011110;
DRAM[35602] = 8'b10011111;
DRAM[35603] = 8'b10011111;
DRAM[35604] = 8'b10011110;
DRAM[35605] = 8'b10011101;
DRAM[35606] = 8'b10011100;
DRAM[35607] = 8'b10011011;
DRAM[35608] = 8'b10011010;
DRAM[35609] = 8'b10011011;
DRAM[35610] = 8'b10011011;
DRAM[35611] = 8'b10011100;
DRAM[35612] = 8'b10011101;
DRAM[35613] = 8'b10011110;
DRAM[35614] = 8'b10011110;
DRAM[35615] = 8'b10011110;
DRAM[35616] = 8'b10100001;
DRAM[35617] = 8'b10100001;
DRAM[35618] = 8'b10100001;
DRAM[35619] = 8'b10100000;
DRAM[35620] = 8'b10100000;
DRAM[35621] = 8'b10100000;
DRAM[35622] = 8'b10100000;
DRAM[35623] = 8'b10100000;
DRAM[35624] = 8'b10100001;
DRAM[35625] = 8'b10100001;
DRAM[35626] = 8'b10100001;
DRAM[35627] = 8'b10100001;
DRAM[35628] = 8'b10100001;
DRAM[35629] = 8'b10100001;
DRAM[35630] = 8'b10100001;
DRAM[35631] = 8'b10100001;
DRAM[35632] = 8'b10011111;
DRAM[35633] = 8'b10011100;
DRAM[35634] = 8'b10011100;
DRAM[35635] = 8'b10011111;
DRAM[35636] = 8'b10100011;
DRAM[35637] = 8'b10101010;
DRAM[35638] = 8'b10111001;
DRAM[35639] = 8'b11000111;
DRAM[35640] = 8'b11000010;
DRAM[35641] = 8'b11000101;
DRAM[35642] = 8'b11001011;
DRAM[35643] = 8'b11011000;
DRAM[35644] = 8'b11101010;
DRAM[35645] = 8'b11110011;
DRAM[35646] = 8'b11101000;
DRAM[35647] = 8'b11010111;
DRAM[35648] = 8'b11001100;
DRAM[35649] = 8'b11000001;
DRAM[35650] = 8'b10110111;
DRAM[35651] = 8'b10110011;
DRAM[35652] = 8'b10101110;
DRAM[35653] = 8'b10100110;
DRAM[35654] = 8'b10011111;
DRAM[35655] = 8'b10011110;
DRAM[35656] = 8'b10100010;
DRAM[35657] = 8'b10100000;
DRAM[35658] = 8'b10011011;
DRAM[35659] = 8'b10010101;
DRAM[35660] = 8'b10010000;
DRAM[35661] = 8'b10001100;
DRAM[35662] = 8'b10001010;
DRAM[35663] = 8'b10001010;
DRAM[35664] = 8'b1111110;
DRAM[35665] = 8'b10001110;
DRAM[35666] = 8'b10011100;
DRAM[35667] = 8'b10011110;
DRAM[35668] = 8'b10011010;
DRAM[35669] = 8'b10011001;
DRAM[35670] = 8'b10011101;
DRAM[35671] = 8'b10100001;
DRAM[35672] = 8'b10011100;
DRAM[35673] = 8'b10100110;
DRAM[35674] = 8'b10110010;
DRAM[35675] = 8'b10111000;
DRAM[35676] = 8'b10110110;
DRAM[35677] = 8'b10110001;
DRAM[35678] = 8'b10101100;
DRAM[35679] = 8'b10101010;
DRAM[35680] = 8'b10100010;
DRAM[35681] = 8'b10100101;
DRAM[35682] = 8'b10100011;
DRAM[35683] = 8'b10011111;
DRAM[35684] = 8'b10011111;
DRAM[35685] = 8'b10100011;
DRAM[35686] = 8'b10100101;
DRAM[35687] = 8'b10100011;
DRAM[35688] = 8'b10101110;
DRAM[35689] = 8'b10101110;
DRAM[35690] = 8'b10100011;
DRAM[35691] = 8'b10011101;
DRAM[35692] = 8'b10100001;
DRAM[35693] = 8'b10011100;
DRAM[35694] = 8'b10100000;
DRAM[35695] = 8'b10110100;
DRAM[35696] = 8'b10111100;
DRAM[35697] = 8'b11001000;
DRAM[35698] = 8'b11001110;
DRAM[35699] = 8'b11000111;
DRAM[35700] = 8'b10111101;
DRAM[35701] = 8'b10111111;
DRAM[35702] = 8'b11001010;
DRAM[35703] = 8'b11010011;
DRAM[35704] = 8'b11100100;
DRAM[35705] = 8'b11100101;
DRAM[35706] = 8'b11100111;
DRAM[35707] = 8'b11101010;
DRAM[35708] = 8'b11101110;
DRAM[35709] = 8'b11110011;
DRAM[35710] = 8'b11110110;
DRAM[35711] = 8'b11111001;
DRAM[35712] = 8'b11111011;
DRAM[35713] = 8'b11111010;
DRAM[35714] = 8'b11111000;
DRAM[35715] = 8'b11110101;
DRAM[35716] = 8'b11110011;
DRAM[35717] = 8'b11110100;
DRAM[35718] = 8'b11110100;
DRAM[35719] = 8'b11110100;
DRAM[35720] = 8'b11110100;
DRAM[35721] = 8'b11110100;
DRAM[35722] = 8'b11110101;
DRAM[35723] = 8'b11110110;
DRAM[35724] = 8'b11110110;
DRAM[35725] = 8'b11110110;
DRAM[35726] = 8'b11110101;
DRAM[35727] = 8'b11110101;
DRAM[35728] = 8'b11110110;
DRAM[35729] = 8'b11110101;
DRAM[35730] = 8'b11110101;
DRAM[35731] = 8'b11110111;
DRAM[35732] = 8'b11111000;
DRAM[35733] = 8'b11111000;
DRAM[35734] = 8'b11110110;
DRAM[35735] = 8'b11110100;
DRAM[35736] = 8'b11110101;
DRAM[35737] = 8'b11110101;
DRAM[35738] = 8'b11110100;
DRAM[35739] = 8'b11110011;
DRAM[35740] = 8'b11110100;
DRAM[35741] = 8'b11110101;
DRAM[35742] = 8'b11110110;
DRAM[35743] = 8'b11110111;
DRAM[35744] = 8'b11111000;
DRAM[35745] = 8'b11110100;
DRAM[35746] = 8'b11110010;
DRAM[35747] = 8'b11110100;
DRAM[35748] = 8'b11110110;
DRAM[35749] = 8'b11110111;
DRAM[35750] = 8'b11111001;
DRAM[35751] = 8'b11111100;
DRAM[35752] = 8'b11101110;
DRAM[35753] = 8'b11101110;
DRAM[35754] = 8'b11101100;
DRAM[35755] = 8'b11100100;
DRAM[35756] = 8'b11010101;
DRAM[35757] = 8'b11001000;
DRAM[35758] = 8'b11000111;
DRAM[35759] = 8'b11001101;
DRAM[35760] = 8'b11010110;
DRAM[35761] = 8'b10110011;
DRAM[35762] = 8'b10100100;
DRAM[35763] = 8'b10111001;
DRAM[35764] = 8'b11001010;
DRAM[35765] = 8'b11000010;
DRAM[35766] = 8'b10111010;
DRAM[35767] = 8'b10111111;
DRAM[35768] = 8'b11000111;
DRAM[35769] = 8'b11000000;
DRAM[35770] = 8'b10110110;
DRAM[35771] = 8'b10110000;
DRAM[35772] = 8'b10101110;
DRAM[35773] = 8'b10101110;
DRAM[35774] = 8'b10101100;
DRAM[35775] = 8'b10101010;
DRAM[35776] = 8'b10100100;
DRAM[35777] = 8'b10010110;
DRAM[35778] = 8'b10001000;
DRAM[35779] = 8'b10000100;
DRAM[35780] = 8'b10001001;
DRAM[35781] = 8'b10010001;
DRAM[35782] = 8'b10011101;
DRAM[35783] = 8'b10100111;
DRAM[35784] = 8'b11000000;
DRAM[35785] = 8'b11001001;
DRAM[35786] = 8'b11010111;
DRAM[35787] = 8'b11100011;
DRAM[35788] = 8'b11101000;
DRAM[35789] = 8'b11011010;
DRAM[35790] = 8'b10111011;
DRAM[35791] = 8'b10011110;
DRAM[35792] = 8'b10001100;
DRAM[35793] = 8'b10010000;
DRAM[35794] = 8'b10010010;
DRAM[35795] = 8'b10001111;
DRAM[35796] = 8'b10001110;
DRAM[35797] = 8'b10010000;
DRAM[35798] = 8'b10001110;
DRAM[35799] = 8'b10001010;
DRAM[35800] = 8'b10001100;
DRAM[35801] = 8'b10001100;
DRAM[35802] = 8'b10001011;
DRAM[35803] = 8'b10001010;
DRAM[35804] = 8'b10001010;
DRAM[35805] = 8'b10001010;
DRAM[35806] = 8'b10001010;
DRAM[35807] = 8'b10001011;
DRAM[35808] = 8'b10001100;
DRAM[35809] = 8'b10001011;
DRAM[35810] = 8'b10001000;
DRAM[35811] = 8'b10000101;
DRAM[35812] = 8'b10000011;
DRAM[35813] = 8'b10000010;
DRAM[35814] = 8'b10000001;
DRAM[35815] = 8'b10000001;
DRAM[35816] = 8'b10000001;
DRAM[35817] = 8'b10000010;
DRAM[35818] = 8'b10000011;
DRAM[35819] = 8'b10000100;
DRAM[35820] = 8'b10000011;
DRAM[35821] = 8'b10000010;
DRAM[35822] = 8'b10000000;
DRAM[35823] = 8'b1111111;
DRAM[35824] = 8'b10000000;
DRAM[35825] = 8'b1111111;
DRAM[35826] = 8'b1111110;
DRAM[35827] = 8'b1111101;
DRAM[35828] = 8'b1111100;
DRAM[35829] = 8'b1111011;
DRAM[35830] = 8'b1111100;
DRAM[35831] = 8'b1111100;
DRAM[35832] = 8'b1111001;
DRAM[35833] = 8'b1111001;
DRAM[35834] = 8'b1111000;
DRAM[35835] = 8'b1111000;
DRAM[35836] = 8'b1111000;
DRAM[35837] = 8'b1110111;
DRAM[35838] = 8'b1110111;
DRAM[35839] = 8'b1110111;
DRAM[35840] = 8'b10010011;
DRAM[35841] = 8'b10010100;
DRAM[35842] = 8'b10010101;
DRAM[35843] = 8'b10010110;
DRAM[35844] = 8'b10011000;
DRAM[35845] = 8'b10011001;
DRAM[35846] = 8'b10011001;
DRAM[35847] = 8'b10011001;
DRAM[35848] = 8'b10011011;
DRAM[35849] = 8'b10011011;
DRAM[35850] = 8'b10011011;
DRAM[35851] = 8'b10011100;
DRAM[35852] = 8'b10011100;
DRAM[35853] = 8'b10011100;
DRAM[35854] = 8'b10011100;
DRAM[35855] = 8'b10011100;
DRAM[35856] = 8'b10011110;
DRAM[35857] = 8'b10011110;
DRAM[35858] = 8'b10011110;
DRAM[35859] = 8'b10011110;
DRAM[35860] = 8'b10011101;
DRAM[35861] = 8'b10011100;
DRAM[35862] = 8'b10011011;
DRAM[35863] = 8'b10011010;
DRAM[35864] = 8'b10011100;
DRAM[35865] = 8'b10011100;
DRAM[35866] = 8'b10011100;
DRAM[35867] = 8'b10011101;
DRAM[35868] = 8'b10011110;
DRAM[35869] = 8'b10011111;
DRAM[35870] = 8'b10011111;
DRAM[35871] = 8'b10100000;
DRAM[35872] = 8'b10100010;
DRAM[35873] = 8'b10100010;
DRAM[35874] = 8'b10100010;
DRAM[35875] = 8'b10100010;
DRAM[35876] = 8'b10100010;
DRAM[35877] = 8'b10100001;
DRAM[35878] = 8'b10100001;
DRAM[35879] = 8'b10100001;
DRAM[35880] = 8'b10100001;
DRAM[35881] = 8'b10100001;
DRAM[35882] = 8'b10100001;
DRAM[35883] = 8'b10100001;
DRAM[35884] = 8'b10100001;
DRAM[35885] = 8'b10100001;
DRAM[35886] = 8'b10100001;
DRAM[35887] = 8'b10100001;
DRAM[35888] = 8'b10100101;
DRAM[35889] = 8'b10100010;
DRAM[35890] = 8'b10100001;
DRAM[35891] = 8'b10100100;
DRAM[35892] = 8'b10101000;
DRAM[35893] = 8'b10101111;
DRAM[35894] = 8'b10111101;
DRAM[35895] = 8'b11001011;
DRAM[35896] = 8'b11011100;
DRAM[35897] = 8'b11100011;
DRAM[35898] = 8'b11100100;
DRAM[35899] = 8'b11100100;
DRAM[35900] = 8'b11101110;
DRAM[35901] = 8'b11111001;
DRAM[35902] = 8'b11110000;
DRAM[35903] = 8'b11011110;
DRAM[35904] = 8'b11001110;
DRAM[35905] = 8'b11000100;
DRAM[35906] = 8'b10111010;
DRAM[35907] = 8'b10110110;
DRAM[35908] = 8'b10110010;
DRAM[35909] = 8'b10101010;
DRAM[35910] = 8'b10100101;
DRAM[35911] = 8'b10100011;
DRAM[35912] = 8'b10100110;
DRAM[35913] = 8'b10100000;
DRAM[35914] = 8'b10011001;
DRAM[35915] = 8'b10010101;
DRAM[35916] = 8'b10010100;
DRAM[35917] = 8'b10010011;
DRAM[35918] = 8'b10001110;
DRAM[35919] = 8'b10001010;
DRAM[35920] = 8'b10001100;
DRAM[35921] = 8'b10011000;
DRAM[35922] = 8'b10100001;
DRAM[35923] = 8'b10100010;
DRAM[35924] = 8'b10100001;
DRAM[35925] = 8'b10100011;
DRAM[35926] = 8'b10100100;
DRAM[35927] = 8'b10100010;
DRAM[35928] = 8'b10100101;
DRAM[35929] = 8'b10101011;
DRAM[35930] = 8'b10110011;
DRAM[35931] = 8'b10110111;
DRAM[35932] = 8'b10110110;
DRAM[35933] = 8'b10110011;
DRAM[35934] = 8'b10110001;
DRAM[35935] = 8'b10110000;
DRAM[35936] = 8'b10100110;
DRAM[35937] = 8'b10100110;
DRAM[35938] = 8'b10100101;
DRAM[35939] = 8'b10100100;
DRAM[35940] = 8'b10101011;
DRAM[35941] = 8'b10110011;
DRAM[35942] = 8'b10110100;
DRAM[35943] = 8'b10101111;
DRAM[35944] = 8'b10110001;
DRAM[35945] = 8'b10101101;
DRAM[35946] = 8'b10101101;
DRAM[35947] = 8'b10100100;
DRAM[35948] = 8'b10010111;
DRAM[35949] = 8'b10100100;
DRAM[35950] = 8'b10111000;
DRAM[35951] = 8'b10111010;
DRAM[35952] = 8'b11001111;
DRAM[35953] = 8'b11000111;
DRAM[35954] = 8'b11000110;
DRAM[35955] = 8'b11001011;
DRAM[35956] = 8'b11001000;
DRAM[35957] = 8'b11000100;
DRAM[35958] = 8'b11001111;
DRAM[35959] = 8'b11100010;
DRAM[35960] = 8'b11100111;
DRAM[35961] = 8'b11100111;
DRAM[35962] = 8'b11101000;
DRAM[35963] = 8'b11101010;
DRAM[35964] = 8'b11101101;
DRAM[35965] = 8'b11110001;
DRAM[35966] = 8'b11110101;
DRAM[35967] = 8'b11110111;
DRAM[35968] = 8'b11110100;
DRAM[35969] = 8'b11110010;
DRAM[35970] = 8'b11101111;
DRAM[35971] = 8'b11101101;
DRAM[35972] = 8'b11101100;
DRAM[35973] = 8'b11101011;
DRAM[35974] = 8'b11101011;
DRAM[35975] = 8'b11101100;
DRAM[35976] = 8'b11110001;
DRAM[35977] = 8'b11110001;
DRAM[35978] = 8'b11110011;
DRAM[35979] = 8'b11110100;
DRAM[35980] = 8'b11110100;
DRAM[35981] = 8'b11110101;
DRAM[35982] = 8'b11110100;
DRAM[35983] = 8'b11110100;
DRAM[35984] = 8'b11101111;
DRAM[35985] = 8'b11101111;
DRAM[35986] = 8'b11110000;
DRAM[35987] = 8'b11110010;
DRAM[35988] = 8'b11110011;
DRAM[35989] = 8'b11110011;
DRAM[35990] = 8'b11110000;
DRAM[35991] = 8'b11101101;
DRAM[35992] = 8'b11101110;
DRAM[35993] = 8'b11110000;
DRAM[35994] = 8'b11110011;
DRAM[35995] = 8'b11110101;
DRAM[35996] = 8'b11110110;
DRAM[35997] = 8'b11110100;
DRAM[35998] = 8'b11110010;
DRAM[35999] = 8'b11110001;
DRAM[36000] = 8'b11110010;
DRAM[36001] = 8'b11101101;
DRAM[36002] = 8'b11101100;
DRAM[36003] = 8'b11110010;
DRAM[36004] = 8'b11110100;
DRAM[36005] = 8'b11110001;
DRAM[36006] = 8'b11101111;
DRAM[36007] = 8'b11110001;
DRAM[36008] = 8'b11101110;
DRAM[36009] = 8'b11101110;
DRAM[36010] = 8'b11110000;
DRAM[36011] = 8'b11101101;
DRAM[36012] = 8'b11011111;
DRAM[36013] = 8'b11001101;
DRAM[36014] = 8'b11000110;
DRAM[36015] = 8'b11001001;
DRAM[36016] = 8'b10111011;
DRAM[36017] = 8'b11001011;
DRAM[36018] = 8'b11000101;
DRAM[36019] = 8'b10101001;
DRAM[36020] = 8'b10100001;
DRAM[36021] = 8'b10111000;
DRAM[36022] = 8'b11001001;
DRAM[36023] = 8'b11000110;
DRAM[36024] = 8'b10110101;
DRAM[36025] = 8'b10110110;
DRAM[36026] = 8'b10111000;
DRAM[36027] = 8'b10111001;
DRAM[36028] = 8'b10110101;
DRAM[36029] = 8'b10101000;
DRAM[36030] = 8'b10011000;
DRAM[36031] = 8'b10001100;
DRAM[36032] = 8'b10011101;
DRAM[36033] = 8'b10010101;
DRAM[36034] = 8'b10010001;
DRAM[36035] = 8'b10010101;
DRAM[36036] = 8'b10011010;
DRAM[36037] = 8'b10011100;
DRAM[36038] = 8'b10011111;
DRAM[36039] = 8'b10100010;
DRAM[36040] = 8'b11000001;
DRAM[36041] = 8'b11001111;
DRAM[36042] = 8'b11011111;
DRAM[36043] = 8'b11100101;
DRAM[36044] = 8'b11100000;
DRAM[36045] = 8'b11001101;
DRAM[36046] = 8'b10110000;
DRAM[36047] = 8'b10011001;
DRAM[36048] = 8'b10001100;
DRAM[36049] = 8'b10010000;
DRAM[36050] = 8'b10010010;
DRAM[36051] = 8'b10001111;
DRAM[36052] = 8'b10001111;
DRAM[36053] = 8'b10010001;
DRAM[36054] = 8'b10001111;
DRAM[36055] = 8'b10001010;
DRAM[36056] = 8'b10001110;
DRAM[36057] = 8'b10001101;
DRAM[36058] = 8'b10001100;
DRAM[36059] = 8'b10001011;
DRAM[36060] = 8'b10001010;
DRAM[36061] = 8'b10001010;
DRAM[36062] = 8'b10001011;
DRAM[36063] = 8'b10001011;
DRAM[36064] = 8'b10001101;
DRAM[36065] = 8'b10001011;
DRAM[36066] = 8'b10001000;
DRAM[36067] = 8'b10000101;
DRAM[36068] = 8'b10000100;
DRAM[36069] = 8'b10000100;
DRAM[36070] = 8'b10000100;
DRAM[36071] = 8'b10000101;
DRAM[36072] = 8'b10000010;
DRAM[36073] = 8'b10000011;
DRAM[36074] = 8'b10000100;
DRAM[36075] = 8'b10000100;
DRAM[36076] = 8'b10000100;
DRAM[36077] = 8'b10000010;
DRAM[36078] = 8'b10000001;
DRAM[36079] = 8'b10000000;
DRAM[36080] = 8'b10000000;
DRAM[36081] = 8'b1111111;
DRAM[36082] = 8'b1111110;
DRAM[36083] = 8'b1111101;
DRAM[36084] = 8'b1111100;
DRAM[36085] = 8'b1111011;
DRAM[36086] = 8'b1111100;
DRAM[36087] = 8'b1111100;
DRAM[36088] = 8'b1111001;
DRAM[36089] = 8'b1111001;
DRAM[36090] = 8'b1111001;
DRAM[36091] = 8'b1111000;
DRAM[36092] = 8'b1111000;
DRAM[36093] = 8'b1111000;
DRAM[36094] = 8'b1110111;
DRAM[36095] = 8'b1110111;
DRAM[36096] = 8'b10010101;
DRAM[36097] = 8'b10010101;
DRAM[36098] = 8'b10010110;
DRAM[36099] = 8'b10010111;
DRAM[36100] = 8'b10011000;
DRAM[36101] = 8'b10011010;
DRAM[36102] = 8'b10011010;
DRAM[36103] = 8'b10011011;
DRAM[36104] = 8'b10011100;
DRAM[36105] = 8'b10011100;
DRAM[36106] = 8'b10011100;
DRAM[36107] = 8'b10011100;
DRAM[36108] = 8'b10011100;
DRAM[36109] = 8'b10011100;
DRAM[36110] = 8'b10011100;
DRAM[36111] = 8'b10011100;
DRAM[36112] = 8'b10011100;
DRAM[36113] = 8'b10011101;
DRAM[36114] = 8'b10011101;
DRAM[36115] = 8'b10011101;
DRAM[36116] = 8'b10011101;
DRAM[36117] = 8'b10011100;
DRAM[36118] = 8'b10011100;
DRAM[36119] = 8'b10011011;
DRAM[36120] = 8'b10011101;
DRAM[36121] = 8'b10011101;
DRAM[36122] = 8'b10011110;
DRAM[36123] = 8'b10011110;
DRAM[36124] = 8'b10011111;
DRAM[36125] = 8'b10100000;
DRAM[36126] = 8'b10100001;
DRAM[36127] = 8'b10100001;
DRAM[36128] = 8'b10100011;
DRAM[36129] = 8'b10100011;
DRAM[36130] = 8'b10100011;
DRAM[36131] = 8'b10100011;
DRAM[36132] = 8'b10100011;
DRAM[36133] = 8'b10100100;
DRAM[36134] = 8'b10100100;
DRAM[36135] = 8'b10100100;
DRAM[36136] = 8'b10100001;
DRAM[36137] = 8'b10100001;
DRAM[36138] = 8'b10100001;
DRAM[36139] = 8'b10100001;
DRAM[36140] = 8'b10100001;
DRAM[36141] = 8'b10100001;
DRAM[36142] = 8'b10100001;
DRAM[36143] = 8'b10100001;
DRAM[36144] = 8'b10100100;
DRAM[36145] = 8'b10100010;
DRAM[36146] = 8'b10100100;
DRAM[36147] = 8'b10101001;
DRAM[36148] = 8'b10101110;
DRAM[36149] = 8'b10110110;
DRAM[36150] = 8'b11000101;
DRAM[36151] = 8'b11010011;
DRAM[36152] = 8'b11100110;
DRAM[36153] = 8'b11110011;
DRAM[36154] = 8'b11111000;
DRAM[36155] = 8'b11110010;
DRAM[36156] = 8'b11110011;
DRAM[36157] = 8'b11111010;
DRAM[36158] = 8'b11110100;
DRAM[36159] = 8'b11100100;
DRAM[36160] = 8'b11010011;
DRAM[36161] = 8'b11001000;
DRAM[36162] = 8'b10111110;
DRAM[36163] = 8'b10111001;
DRAM[36164] = 8'b10110101;
DRAM[36165] = 8'b10101110;
DRAM[36166] = 8'b10101010;
DRAM[36167] = 8'b10101001;
DRAM[36168] = 8'b10100100;
DRAM[36169] = 8'b10011101;
DRAM[36170] = 8'b10010101;
DRAM[36171] = 8'b10010010;
DRAM[36172] = 8'b10010100;
DRAM[36173] = 8'b10010100;
DRAM[36174] = 8'b10001111;
DRAM[36175] = 8'b10001001;
DRAM[36176] = 8'b10010110;
DRAM[36177] = 8'b10011110;
DRAM[36178] = 8'b10100011;
DRAM[36179] = 8'b10100010;
DRAM[36180] = 8'b10100100;
DRAM[36181] = 8'b10101010;
DRAM[36182] = 8'b10101010;
DRAM[36183] = 8'b10100100;
DRAM[36184] = 8'b10101111;
DRAM[36185] = 8'b10101110;
DRAM[36186] = 8'b10101100;
DRAM[36187] = 8'b10101011;
DRAM[36188] = 8'b10101110;
DRAM[36189] = 8'b10110001;
DRAM[36190] = 8'b10110101;
DRAM[36191] = 8'b10111000;
DRAM[36192] = 8'b11000001;
DRAM[36193] = 8'b10111011;
DRAM[36194] = 8'b10110110;
DRAM[36195] = 8'b10110100;
DRAM[36196] = 8'b10110100;
DRAM[36197] = 8'b10110001;
DRAM[36198] = 8'b10101011;
DRAM[36199] = 8'b10100110;
DRAM[36200] = 8'b10010111;
DRAM[36201] = 8'b10011001;
DRAM[36202] = 8'b10100101;
DRAM[36203] = 8'b10100010;
DRAM[36204] = 8'b10011011;
DRAM[36205] = 8'b10110011;
DRAM[36206] = 8'b11001000;
DRAM[36207] = 8'b10111110;
DRAM[36208] = 8'b11001100;
DRAM[36209] = 8'b10111011;
DRAM[36210] = 8'b10111010;
DRAM[36211] = 8'b11001001;
DRAM[36212] = 8'b11001111;
DRAM[36213] = 8'b11001010;
DRAM[36214] = 8'b11010100;
DRAM[36215] = 8'b11101001;
DRAM[36216] = 8'b11100100;
DRAM[36217] = 8'b11100110;
DRAM[36218] = 8'b11101010;
DRAM[36219] = 8'b11101110;
DRAM[36220] = 8'b11110001;
DRAM[36221] = 8'b11110001;
DRAM[36222] = 8'b11110001;
DRAM[36223] = 8'b11110000;
DRAM[36224] = 8'b11110001;
DRAM[36225] = 8'b11101110;
DRAM[36226] = 8'b11101100;
DRAM[36227] = 8'b11101101;
DRAM[36228] = 8'b11101100;
DRAM[36229] = 8'b11101000;
DRAM[36230] = 8'b11101000;
DRAM[36231] = 8'b11101010;
DRAM[36232] = 8'b11110000;
DRAM[36233] = 8'b11110001;
DRAM[36234] = 8'b11110001;
DRAM[36235] = 8'b11110010;
DRAM[36236] = 8'b11110010;
DRAM[36237] = 8'b11110001;
DRAM[36238] = 8'b11110001;
DRAM[36239] = 8'b11110000;
DRAM[36240] = 8'b11101011;
DRAM[36241] = 8'b11101001;
DRAM[36242] = 8'b11101000;
DRAM[36243] = 8'b11101000;
DRAM[36244] = 8'b11101010;
DRAM[36245] = 8'b11101010;
DRAM[36246] = 8'b11101010;
DRAM[36247] = 8'b11101000;
DRAM[36248] = 8'b11100111;
DRAM[36249] = 8'b11101011;
DRAM[36250] = 8'b11110000;
DRAM[36251] = 8'b11110101;
DRAM[36252] = 8'b11110111;
DRAM[36253] = 8'b11110110;
DRAM[36254] = 8'b11110011;
DRAM[36255] = 8'b11110001;
DRAM[36256] = 8'b11110001;
DRAM[36257] = 8'b11101010;
DRAM[36258] = 8'b11101010;
DRAM[36259] = 8'b11110010;
DRAM[36260] = 8'b11110101;
DRAM[36261] = 8'b11101111;
DRAM[36262] = 8'b11101010;
DRAM[36263] = 8'b11101011;
DRAM[36264] = 8'b11101110;
DRAM[36265] = 8'b11101110;
DRAM[36266] = 8'b11101111;
DRAM[36267] = 8'b11101111;
DRAM[36268] = 8'b11100111;
DRAM[36269] = 8'b11010110;
DRAM[36270] = 8'b11000110;
DRAM[36271] = 8'b10111110;
DRAM[36272] = 8'b10100101;
DRAM[36273] = 8'b11000100;
DRAM[36274] = 8'b11010001;
DRAM[36275] = 8'b10111011;
DRAM[36276] = 8'b10100100;
DRAM[36277] = 8'b10100110;
DRAM[36278] = 8'b10110100;
DRAM[36279] = 8'b10111011;
DRAM[36280] = 8'b10111110;
DRAM[36281] = 8'b10110100;
DRAM[36282] = 8'b10101001;
DRAM[36283] = 8'b10100011;
DRAM[36284] = 8'b10100101;
DRAM[36285] = 8'b10101011;
DRAM[36286] = 8'b10110000;
DRAM[36287] = 8'b10110010;
DRAM[36288] = 8'b10011010;
DRAM[36289] = 8'b10010100;
DRAM[36290] = 8'b10010001;
DRAM[36291] = 8'b10010101;
DRAM[36292] = 8'b10011100;
DRAM[36293] = 8'b10100001;
DRAM[36294] = 8'b10101010;
DRAM[36295] = 8'b10110001;
DRAM[36296] = 8'b10110011;
DRAM[36297] = 8'b11001111;
DRAM[36298] = 8'b11101001;
DRAM[36299] = 8'b11101011;
DRAM[36300] = 8'b11011000;
DRAM[36301] = 8'b11000011;
DRAM[36302] = 8'b10110011;
DRAM[36303] = 8'b10101011;
DRAM[36304] = 8'b10011001;
DRAM[36305] = 8'b10010110;
DRAM[36306] = 8'b10010011;
DRAM[36307] = 8'b10010010;
DRAM[36308] = 8'b10010010;
DRAM[36309] = 8'b10010010;
DRAM[36310] = 8'b10010000;
DRAM[36311] = 8'b10001111;
DRAM[36312] = 8'b10001111;
DRAM[36313] = 8'b10001110;
DRAM[36314] = 8'b10001101;
DRAM[36315] = 8'b10001100;
DRAM[36316] = 8'b10001011;
DRAM[36317] = 8'b10001011;
DRAM[36318] = 8'b10001011;
DRAM[36319] = 8'b10001011;
DRAM[36320] = 8'b10001011;
DRAM[36321] = 8'b10001010;
DRAM[36322] = 8'b10001000;
DRAM[36323] = 8'b10000110;
DRAM[36324] = 8'b10000101;
DRAM[36325] = 8'b10000101;
DRAM[36326] = 8'b10000110;
DRAM[36327] = 8'b10000110;
DRAM[36328] = 8'b10000010;
DRAM[36329] = 8'b10000011;
DRAM[36330] = 8'b10000011;
DRAM[36331] = 8'b10000011;
DRAM[36332] = 8'b10000011;
DRAM[36333] = 8'b10000010;
DRAM[36334] = 8'b10000001;
DRAM[36335] = 8'b10000000;
DRAM[36336] = 8'b10000000;
DRAM[36337] = 8'b1111111;
DRAM[36338] = 8'b1111110;
DRAM[36339] = 8'b1111101;
DRAM[36340] = 8'b1111100;
DRAM[36341] = 8'b1111011;
DRAM[36342] = 8'b1111100;
DRAM[36343] = 8'b1111100;
DRAM[36344] = 8'b1111010;
DRAM[36345] = 8'b1111001;
DRAM[36346] = 8'b1111001;
DRAM[36347] = 8'b1111001;
DRAM[36348] = 8'b1111000;
DRAM[36349] = 8'b1111000;
DRAM[36350] = 8'b1111000;
DRAM[36351] = 8'b1111000;
DRAM[36352] = 8'b10010110;
DRAM[36353] = 8'b10010110;
DRAM[36354] = 8'b10010111;
DRAM[36355] = 8'b10011000;
DRAM[36356] = 8'b10011001;
DRAM[36357] = 8'b10011010;
DRAM[36358] = 8'b10011100;
DRAM[36359] = 8'b10011100;
DRAM[36360] = 8'b10011100;
DRAM[36361] = 8'b10011100;
DRAM[36362] = 8'b10011100;
DRAM[36363] = 8'b10011100;
DRAM[36364] = 8'b10011100;
DRAM[36365] = 8'b10011100;
DRAM[36366] = 8'b10011100;
DRAM[36367] = 8'b10011100;
DRAM[36368] = 8'b10011100;
DRAM[36369] = 8'b10011100;
DRAM[36370] = 8'b10011101;
DRAM[36371] = 8'b10011110;
DRAM[36372] = 8'b10011110;
DRAM[36373] = 8'b10011110;
DRAM[36374] = 8'b10011101;
DRAM[36375] = 8'b10011101;
DRAM[36376] = 8'b10011110;
DRAM[36377] = 8'b10011110;
DRAM[36378] = 8'b10011110;
DRAM[36379] = 8'b10011111;
DRAM[36380] = 8'b10100000;
DRAM[36381] = 8'b10100001;
DRAM[36382] = 8'b10100001;
DRAM[36383] = 8'b10100010;
DRAM[36384] = 8'b10100011;
DRAM[36385] = 8'b10100011;
DRAM[36386] = 8'b10100100;
DRAM[36387] = 8'b10100100;
DRAM[36388] = 8'b10100101;
DRAM[36389] = 8'b10100101;
DRAM[36390] = 8'b10100110;
DRAM[36391] = 8'b10100110;
DRAM[36392] = 8'b10100011;
DRAM[36393] = 8'b10100011;
DRAM[36394] = 8'b10100011;
DRAM[36395] = 8'b10100011;
DRAM[36396] = 8'b10100011;
DRAM[36397] = 8'b10100011;
DRAM[36398] = 8'b10100011;
DRAM[36399] = 8'b10100011;
DRAM[36400] = 8'b10100010;
DRAM[36401] = 8'b10100001;
DRAM[36402] = 8'b10100011;
DRAM[36403] = 8'b10101000;
DRAM[36404] = 8'b10101101;
DRAM[36405] = 8'b10110100;
DRAM[36406] = 8'b11000001;
DRAM[36407] = 8'b11001101;
DRAM[36408] = 8'b11010110;
DRAM[36409] = 8'b11101010;
DRAM[36410] = 8'b11111010;
DRAM[36411] = 8'b11111100;
DRAM[36412] = 8'b11111100;
DRAM[36413] = 8'b11111110;
DRAM[36414] = 8'b11110110;
DRAM[36415] = 8'b11101000;
DRAM[36416] = 8'b11011010;
DRAM[36417] = 8'b11001110;
DRAM[36418] = 8'b11000010;
DRAM[36419] = 8'b10111100;
DRAM[36420] = 8'b10110111;
DRAM[36421] = 8'b10110000;
DRAM[36422] = 8'b10101100;
DRAM[36423] = 8'b10101100;
DRAM[36424] = 8'b10100011;
DRAM[36425] = 8'b10011111;
DRAM[36426] = 8'b10011010;
DRAM[36427] = 8'b10010111;
DRAM[36428] = 8'b10010111;
DRAM[36429] = 8'b10010110;
DRAM[36430] = 8'b10010011;
DRAM[36431] = 8'b10010001;
DRAM[36432] = 8'b10001011;
DRAM[36433] = 8'b10010101;
DRAM[36434] = 8'b10011000;
DRAM[36435] = 8'b10010100;
DRAM[36436] = 8'b10010110;
DRAM[36437] = 8'b10011111;
DRAM[36438] = 8'b10100001;
DRAM[36439] = 8'b10011100;
DRAM[36440] = 8'b10101101;
DRAM[36441] = 8'b10101001;
DRAM[36442] = 8'b10100110;
DRAM[36443] = 8'b10100111;
DRAM[36444] = 8'b10101110;
DRAM[36445] = 8'b10110100;
DRAM[36446] = 8'b10110111;
DRAM[36447] = 8'b10110111;
DRAM[36448] = 8'b10111000;
DRAM[36449] = 8'b10110010;
DRAM[36450] = 8'b10110011;
DRAM[36451] = 8'b10111000;
DRAM[36452] = 8'b10110111;
DRAM[36453] = 8'b10101110;
DRAM[36454] = 8'b10101100;
DRAM[36455] = 8'b10101111;
DRAM[36456] = 8'b10110011;
DRAM[36457] = 8'b10111100;
DRAM[36458] = 8'b10110011;
DRAM[36459] = 8'b10101011;
DRAM[36460] = 8'b10110101;
DRAM[36461] = 8'b10111101;
DRAM[36462] = 8'b10111001;
DRAM[36463] = 8'b10110110;
DRAM[36464] = 8'b10111100;
DRAM[36465] = 8'b10110101;
DRAM[36466] = 8'b10111001;
DRAM[36467] = 8'b11000111;
DRAM[36468] = 8'b11001111;
DRAM[36469] = 8'b11001111;
DRAM[36470] = 8'b11010111;
DRAM[36471] = 8'b11100100;
DRAM[36472] = 8'b11100101;
DRAM[36473] = 8'b11100111;
DRAM[36474] = 8'b11101001;
DRAM[36475] = 8'b11101011;
DRAM[36476] = 8'b11101101;
DRAM[36477] = 8'b11101110;
DRAM[36478] = 8'b11101110;
DRAM[36479] = 8'b11101110;
DRAM[36480] = 8'b11110001;
DRAM[36481] = 8'b11101101;
DRAM[36482] = 8'b11101101;
DRAM[36483] = 8'b11110000;
DRAM[36484] = 8'b11101111;
DRAM[36485] = 8'b11101010;
DRAM[36486] = 8'b11101000;
DRAM[36487] = 8'b11101011;
DRAM[36488] = 8'b11101111;
DRAM[36489] = 8'b11101110;
DRAM[36490] = 8'b11101101;
DRAM[36491] = 8'b11101100;
DRAM[36492] = 8'b11101010;
DRAM[36493] = 8'b11100111;
DRAM[36494] = 8'b11100101;
DRAM[36495] = 8'b11100100;
DRAM[36496] = 8'b11011101;
DRAM[36497] = 8'b11010111;
DRAM[36498] = 8'b11010001;
DRAM[36499] = 8'b11001110;
DRAM[36500] = 8'b11001111;
DRAM[36501] = 8'b11010100;
DRAM[36502] = 8'b11011000;
DRAM[36503] = 8'b11011010;
DRAM[36504] = 8'b11011001;
DRAM[36505] = 8'b11011101;
DRAM[36506] = 8'b11100011;
DRAM[36507] = 8'b11101010;
DRAM[36508] = 8'b11101110;
DRAM[36509] = 8'b11110000;
DRAM[36510] = 8'b11110000;
DRAM[36511] = 8'b11101111;
DRAM[36512] = 8'b11100101;
DRAM[36513] = 8'b11011101;
DRAM[36514] = 8'b11011110;
DRAM[36515] = 8'b11101011;
DRAM[36516] = 8'b11110010;
DRAM[36517] = 8'b11101110;
DRAM[36518] = 8'b11101100;
DRAM[36519] = 8'b11101111;
DRAM[36520] = 8'b11110001;
DRAM[36521] = 8'b11101101;
DRAM[36522] = 8'b11101010;
DRAM[36523] = 8'b11101010;
DRAM[36524] = 8'b11101001;
DRAM[36525] = 8'b11011111;
DRAM[36526] = 8'b11001000;
DRAM[36527] = 8'b10110010;
DRAM[36528] = 8'b11000000;
DRAM[36529] = 8'b10101001;
DRAM[36530] = 8'b10100101;
DRAM[36531] = 8'b11000000;
DRAM[36532] = 8'b11010010;
DRAM[36533] = 8'b11000111;
DRAM[36534] = 8'b10110001;
DRAM[36535] = 8'b10100110;
DRAM[36536] = 8'b11000010;
DRAM[36537] = 8'b11000011;
DRAM[36538] = 8'b11000100;
DRAM[36539] = 8'b11000101;
DRAM[36540] = 8'b11000001;
DRAM[36541] = 8'b10110110;
DRAM[36542] = 8'b10100110;
DRAM[36543] = 8'b10011010;
DRAM[36544] = 8'b10011011;
DRAM[36545] = 8'b10010101;
DRAM[36546] = 8'b10010000;
DRAM[36547] = 8'b10010001;
DRAM[36548] = 8'b10010110;
DRAM[36549] = 8'b10100000;
DRAM[36550] = 8'b10110000;
DRAM[36551] = 8'b10111110;
DRAM[36552] = 8'b10111111;
DRAM[36553] = 8'b11011001;
DRAM[36554] = 8'b11110011;
DRAM[36555] = 8'b11110111;
DRAM[36556] = 8'b11101010;
DRAM[36557] = 8'b11011001;
DRAM[36558] = 8'b11001100;
DRAM[36559] = 8'b11000101;
DRAM[36560] = 8'b10101001;
DRAM[36561] = 8'b10011011;
DRAM[36562] = 8'b10010001;
DRAM[36563] = 8'b10010010;
DRAM[36564] = 8'b10010011;
DRAM[36565] = 8'b10001111;
DRAM[36566] = 8'b10001110;
DRAM[36567] = 8'b10010001;
DRAM[36568] = 8'b10010000;
DRAM[36569] = 8'b10001111;
DRAM[36570] = 8'b10001110;
DRAM[36571] = 8'b10001100;
DRAM[36572] = 8'b10001011;
DRAM[36573] = 8'b10001011;
DRAM[36574] = 8'b10001011;
DRAM[36575] = 8'b10001011;
DRAM[36576] = 8'b10001010;
DRAM[36577] = 8'b10001001;
DRAM[36578] = 8'b10001000;
DRAM[36579] = 8'b10000110;
DRAM[36580] = 8'b10000101;
DRAM[36581] = 8'b10000100;
DRAM[36582] = 8'b10000100;
DRAM[36583] = 8'b10000100;
DRAM[36584] = 8'b10000011;
DRAM[36585] = 8'b10000011;
DRAM[36586] = 8'b10000010;
DRAM[36587] = 8'b10000001;
DRAM[36588] = 8'b10000001;
DRAM[36589] = 8'b10000001;
DRAM[36590] = 8'b10000001;
DRAM[36591] = 8'b10000001;
DRAM[36592] = 8'b10000000;
DRAM[36593] = 8'b1111111;
DRAM[36594] = 8'b1111110;
DRAM[36595] = 8'b1111101;
DRAM[36596] = 8'b1111100;
DRAM[36597] = 8'b1111011;
DRAM[36598] = 8'b1111100;
DRAM[36599] = 8'b1111100;
DRAM[36600] = 8'b1111010;
DRAM[36601] = 8'b1111010;
DRAM[36602] = 8'b1111001;
DRAM[36603] = 8'b1111001;
DRAM[36604] = 8'b1111001;
DRAM[36605] = 8'b1111000;
DRAM[36606] = 8'b1111000;
DRAM[36607] = 8'b1111000;
DRAM[36608] = 8'b10010111;
DRAM[36609] = 8'b10010111;
DRAM[36610] = 8'b10010111;
DRAM[36611] = 8'b10011000;
DRAM[36612] = 8'b10011001;
DRAM[36613] = 8'b10011011;
DRAM[36614] = 8'b10011100;
DRAM[36615] = 8'b10011101;
DRAM[36616] = 8'b10011100;
DRAM[36617] = 8'b10011100;
DRAM[36618] = 8'b10011100;
DRAM[36619] = 8'b10011100;
DRAM[36620] = 8'b10011100;
DRAM[36621] = 8'b10011100;
DRAM[36622] = 8'b10011100;
DRAM[36623] = 8'b10011100;
DRAM[36624] = 8'b10011100;
DRAM[36625] = 8'b10011100;
DRAM[36626] = 8'b10011101;
DRAM[36627] = 8'b10011110;
DRAM[36628] = 8'b10011111;
DRAM[36629] = 8'b10011111;
DRAM[36630] = 8'b10011111;
DRAM[36631] = 8'b10011111;
DRAM[36632] = 8'b10011110;
DRAM[36633] = 8'b10011110;
DRAM[36634] = 8'b10011111;
DRAM[36635] = 8'b10100000;
DRAM[36636] = 8'b10100001;
DRAM[36637] = 8'b10100001;
DRAM[36638] = 8'b10100010;
DRAM[36639] = 8'b10100010;
DRAM[36640] = 8'b10100011;
DRAM[36641] = 8'b10100011;
DRAM[36642] = 8'b10100100;
DRAM[36643] = 8'b10100101;
DRAM[36644] = 8'b10100110;
DRAM[36645] = 8'b10100111;
DRAM[36646] = 8'b10100111;
DRAM[36647] = 8'b10101000;
DRAM[36648] = 8'b10100100;
DRAM[36649] = 8'b10100100;
DRAM[36650] = 8'b10100100;
DRAM[36651] = 8'b10100100;
DRAM[36652] = 8'b10100100;
DRAM[36653] = 8'b10100100;
DRAM[36654] = 8'b10100100;
DRAM[36655] = 8'b10100100;
DRAM[36656] = 8'b10101010;
DRAM[36657] = 8'b10100111;
DRAM[36658] = 8'b10100110;
DRAM[36659] = 8'b10100110;
DRAM[36660] = 8'b10100101;
DRAM[36661] = 8'b10100110;
DRAM[36662] = 8'b10101110;
DRAM[36663] = 8'b10111000;
DRAM[36664] = 8'b11001100;
DRAM[36665] = 8'b11011110;
DRAM[36666] = 8'b11101110;
DRAM[36667] = 8'b11110011;
DRAM[36668] = 8'b11110111;
DRAM[36669] = 8'b11111101;
DRAM[36670] = 8'b11111100;
DRAM[36671] = 8'b11110101;
DRAM[36672] = 8'b11011111;
DRAM[36673] = 8'b11010010;
DRAM[36674] = 8'b11000101;
DRAM[36675] = 8'b10111101;
DRAM[36676] = 8'b10110111;
DRAM[36677] = 8'b10110000;
DRAM[36678] = 8'b10101100;
DRAM[36679] = 8'b10101100;
DRAM[36680] = 8'b10100110;
DRAM[36681] = 8'b10100110;
DRAM[36682] = 8'b10100100;
DRAM[36683] = 8'b10100000;
DRAM[36684] = 8'b10011100;
DRAM[36685] = 8'b10011010;
DRAM[36686] = 8'b10011011;
DRAM[36687] = 8'b10011101;
DRAM[36688] = 8'b10010100;
DRAM[36689] = 8'b10100000;
DRAM[36690] = 8'b10100100;
DRAM[36691] = 8'b10011110;
DRAM[36692] = 8'b10011101;
DRAM[36693] = 8'b10100111;
DRAM[36694] = 8'b10101101;
DRAM[36695] = 8'b10101010;
DRAM[36696] = 8'b10101001;
DRAM[36697] = 8'b10100111;
DRAM[36698] = 8'b10101001;
DRAM[36699] = 8'b10110001;
DRAM[36700] = 8'b10111011;
DRAM[36701] = 8'b10111111;
DRAM[36702] = 8'b10111011;
DRAM[36703] = 8'b10110101;
DRAM[36704] = 8'b10111101;
DRAM[36705] = 8'b10110111;
DRAM[36706] = 8'b10111001;
DRAM[36707] = 8'b10111101;
DRAM[36708] = 8'b10110010;
DRAM[36709] = 8'b10011111;
DRAM[36710] = 8'b10011011;
DRAM[36711] = 8'b10100100;
DRAM[36712] = 8'b10110111;
DRAM[36713] = 8'b11000100;
DRAM[36714] = 8'b10100110;
DRAM[36715] = 8'b10011100;
DRAM[36716] = 8'b11000010;
DRAM[36717] = 8'b10111111;
DRAM[36718] = 8'b10101001;
DRAM[36719] = 8'b10111011;
DRAM[36720] = 8'b10110100;
DRAM[36721] = 8'b10111011;
DRAM[36722] = 8'b11000100;
DRAM[36723] = 8'b11001100;
DRAM[36724] = 8'b11010001;
DRAM[36725] = 8'b11010111;
DRAM[36726] = 8'b11011100;
DRAM[36727] = 8'b11011111;
DRAM[36728] = 8'b11101101;
DRAM[36729] = 8'b11101001;
DRAM[36730] = 8'b11100101;
DRAM[36731] = 8'b11100011;
DRAM[36732] = 8'b11100100;
DRAM[36733] = 8'b11101001;
DRAM[36734] = 8'b11101111;
DRAM[36735] = 8'b11110100;
DRAM[36736] = 8'b11101100;
DRAM[36737] = 8'b11101000;
DRAM[36738] = 8'b11101001;
DRAM[36739] = 8'b11101110;
DRAM[36740] = 8'b11101101;
DRAM[36741] = 8'b11100111;
DRAM[36742] = 8'b11100101;
DRAM[36743] = 8'b11101000;
DRAM[36744] = 8'b11101011;
DRAM[36745] = 8'b11101010;
DRAM[36746] = 8'b11101000;
DRAM[36747] = 8'b11100101;
DRAM[36748] = 8'b11100001;
DRAM[36749] = 8'b11011101;
DRAM[36750] = 8'b11011001;
DRAM[36751] = 8'b11010111;
DRAM[36752] = 8'b11001000;
DRAM[36753] = 8'b11000000;
DRAM[36754] = 8'b10110101;
DRAM[36755] = 8'b10101110;
DRAM[36756] = 8'b10110000;
DRAM[36757] = 8'b10110111;
DRAM[36758] = 8'b11000000;
DRAM[36759] = 8'b11000110;
DRAM[36760] = 8'b11000110;
DRAM[36761] = 8'b11001010;
DRAM[36762] = 8'b11010000;
DRAM[36763] = 8'b11010111;
DRAM[36764] = 8'b11011110;
DRAM[36765] = 8'b11100011;
DRAM[36766] = 8'b11100110;
DRAM[36767] = 8'b11100111;
DRAM[36768] = 8'b11010001;
DRAM[36769] = 8'b11001001;
DRAM[36770] = 8'b11001100;
DRAM[36771] = 8'b11011100;
DRAM[36772] = 8'b11101000;
DRAM[36773] = 8'b11101001;
DRAM[36774] = 8'b11101011;
DRAM[36775] = 8'b11110001;
DRAM[36776] = 8'b11110111;
DRAM[36777] = 8'b11110001;
DRAM[36778] = 8'b11101001;
DRAM[36779] = 8'b11101000;
DRAM[36780] = 8'b11101101;
DRAM[36781] = 8'b11101000;
DRAM[36782] = 8'b11001101;
DRAM[36783] = 8'b10101111;
DRAM[36784] = 8'b10110001;
DRAM[36785] = 8'b10110101;
DRAM[36786] = 8'b10111000;
DRAM[36787] = 8'b10111010;
DRAM[36788] = 8'b10111101;
DRAM[36789] = 8'b11000010;
DRAM[36790] = 8'b11001010;
DRAM[36791] = 8'b11010000;
DRAM[36792] = 8'b11001010;
DRAM[36793] = 8'b11001001;
DRAM[36794] = 8'b11000111;
DRAM[36795] = 8'b11000101;
DRAM[36796] = 8'b10111111;
DRAM[36797] = 8'b10110011;
DRAM[36798] = 8'b10100011;
DRAM[36799] = 8'b10011000;
DRAM[36800] = 8'b10010000;
DRAM[36801] = 8'b10010001;
DRAM[36802] = 8'b10010110;
DRAM[36803] = 8'b10011101;
DRAM[36804] = 8'b10100000;
DRAM[36805] = 8'b10100010;
DRAM[36806] = 8'b10101001;
DRAM[36807] = 8'b10110010;
DRAM[36808] = 8'b11000111;
DRAM[36809] = 8'b11010100;
DRAM[36810] = 8'b11100011;
DRAM[36811] = 8'b11101101;
DRAM[36812] = 8'b11110000;
DRAM[36813] = 8'b11100111;
DRAM[36814] = 8'b11010010;
DRAM[36815] = 8'b10111110;
DRAM[36816] = 8'b10110010;
DRAM[36817] = 8'b10011100;
DRAM[36818] = 8'b10001101;
DRAM[36819] = 8'b10010000;
DRAM[36820] = 8'b10010001;
DRAM[36821] = 8'b10001011;
DRAM[36822] = 8'b10001010;
DRAM[36823] = 8'b10010000;
DRAM[36824] = 8'b10010000;
DRAM[36825] = 8'b10010000;
DRAM[36826] = 8'b10001110;
DRAM[36827] = 8'b10001101;
DRAM[36828] = 8'b10001100;
DRAM[36829] = 8'b10001011;
DRAM[36830] = 8'b10001011;
DRAM[36831] = 8'b10001011;
DRAM[36832] = 8'b10001010;
DRAM[36833] = 8'b10001001;
DRAM[36834] = 8'b10001000;
DRAM[36835] = 8'b10000110;
DRAM[36836] = 8'b10000100;
DRAM[36837] = 8'b10000010;
DRAM[36838] = 8'b10000001;
DRAM[36839] = 8'b10000000;
DRAM[36840] = 8'b10000100;
DRAM[36841] = 8'b10000010;
DRAM[36842] = 8'b10000001;
DRAM[36843] = 8'b1111111;
DRAM[36844] = 8'b1111111;
DRAM[36845] = 8'b10000000;
DRAM[36846] = 8'b10000001;
DRAM[36847] = 8'b10000010;
DRAM[36848] = 8'b10000000;
DRAM[36849] = 8'b1111111;
DRAM[36850] = 8'b1111110;
DRAM[36851] = 8'b1111101;
DRAM[36852] = 8'b1111100;
DRAM[36853] = 8'b1111011;
DRAM[36854] = 8'b1111100;
DRAM[36855] = 8'b1111100;
DRAM[36856] = 8'b1111010;
DRAM[36857] = 8'b1111010;
DRAM[36858] = 8'b1111010;
DRAM[36859] = 8'b1111001;
DRAM[36860] = 8'b1111001;
DRAM[36861] = 8'b1111000;
DRAM[36862] = 8'b1111000;
DRAM[36863] = 8'b1111000;
DRAM[36864] = 8'b10011000;
DRAM[36865] = 8'b10011000;
DRAM[36866] = 8'b10011001;
DRAM[36867] = 8'b10011010;
DRAM[36868] = 8'b10011010;
DRAM[36869] = 8'b10011011;
DRAM[36870] = 8'b10011100;
DRAM[36871] = 8'b10011100;
DRAM[36872] = 8'b10011101;
DRAM[36873] = 8'b10011101;
DRAM[36874] = 8'b10011110;
DRAM[36875] = 8'b10011110;
DRAM[36876] = 8'b10011110;
DRAM[36877] = 8'b10011110;
DRAM[36878] = 8'b10011111;
DRAM[36879] = 8'b10011111;
DRAM[36880] = 8'b10100000;
DRAM[36881] = 8'b10011111;
DRAM[36882] = 8'b10011111;
DRAM[36883] = 8'b10011111;
DRAM[36884] = 8'b10011111;
DRAM[36885] = 8'b10100000;
DRAM[36886] = 8'b10100001;
DRAM[36887] = 8'b10100010;
DRAM[36888] = 8'b10011111;
DRAM[36889] = 8'b10011111;
DRAM[36890] = 8'b10011111;
DRAM[36891] = 8'b10100000;
DRAM[36892] = 8'b10100001;
DRAM[36893] = 8'b10100010;
DRAM[36894] = 8'b10100011;
DRAM[36895] = 8'b10100100;
DRAM[36896] = 8'b10100101;
DRAM[36897] = 8'b10100110;
DRAM[36898] = 8'b10100111;
DRAM[36899] = 8'b10101000;
DRAM[36900] = 8'b10101000;
DRAM[36901] = 8'b10101000;
DRAM[36902] = 8'b10101000;
DRAM[36903] = 8'b10101000;
DRAM[36904] = 8'b10100101;
DRAM[36905] = 8'b10100100;
DRAM[36906] = 8'b10100100;
DRAM[36907] = 8'b10100011;
DRAM[36908] = 8'b10100011;
DRAM[36909] = 8'b10100100;
DRAM[36910] = 8'b10100100;
DRAM[36911] = 8'b10100101;
DRAM[36912] = 8'b10100000;
DRAM[36913] = 8'b10100010;
DRAM[36914] = 8'b10100011;
DRAM[36915] = 8'b10100001;
DRAM[36916] = 8'b10100001;
DRAM[36917] = 8'b10100111;
DRAM[36918] = 8'b10110001;
DRAM[36919] = 8'b10111010;
DRAM[36920] = 8'b10111011;
DRAM[36921] = 8'b11010000;
DRAM[36922] = 8'b11100111;
DRAM[36923] = 8'b11110110;
DRAM[36924] = 8'b11111011;
DRAM[36925] = 8'b11111100;
DRAM[36926] = 8'b11111000;
DRAM[36927] = 8'b11110011;
DRAM[36928] = 8'b11011111;
DRAM[36929] = 8'b11010110;
DRAM[36930] = 8'b11001010;
DRAM[36931] = 8'b11000001;
DRAM[36932] = 8'b10111010;
DRAM[36933] = 8'b10110101;
DRAM[36934] = 8'b10101111;
DRAM[36935] = 8'b10101011;
DRAM[36936] = 8'b10110000;
DRAM[36937] = 8'b10101100;
DRAM[36938] = 8'b10101001;
DRAM[36939] = 8'b10101000;
DRAM[36940] = 8'b10101000;
DRAM[36941] = 8'b10100011;
DRAM[36942] = 8'b10011000;
DRAM[36943] = 8'b10010000;
DRAM[36944] = 8'b10001100;
DRAM[36945] = 8'b10100000;
DRAM[36946] = 8'b10100010;
DRAM[36947] = 8'b10011011;
DRAM[36948] = 8'b10010111;
DRAM[36949] = 8'b10001010;
DRAM[36950] = 8'b10010001;
DRAM[36951] = 8'b10110001;
DRAM[36952] = 8'b10110100;
DRAM[36953] = 8'b10110100;
DRAM[36954] = 8'b10110011;
DRAM[36955] = 8'b10110010;
DRAM[36956] = 8'b10110001;
DRAM[36957] = 8'b10110101;
DRAM[36958] = 8'b10111100;
DRAM[36959] = 8'b11000010;
DRAM[36960] = 8'b10111011;
DRAM[36961] = 8'b10110100;
DRAM[36962] = 8'b10101100;
DRAM[36963] = 8'b10101011;
DRAM[36964] = 8'b10110001;
DRAM[36965] = 8'b10111001;
DRAM[36966] = 8'b10111101;
DRAM[36967] = 8'b10111110;
DRAM[36968] = 8'b10101111;
DRAM[36969] = 8'b10010011;
DRAM[36970] = 8'b10010100;
DRAM[36971] = 8'b10111001;
DRAM[36972] = 8'b11001011;
DRAM[36973] = 8'b10111011;
DRAM[36974] = 8'b10110101;
DRAM[36975] = 8'b11000010;
DRAM[36976] = 8'b10110010;
DRAM[36977] = 8'b11000001;
DRAM[36978] = 8'b11001010;
DRAM[36979] = 8'b11001001;
DRAM[36980] = 8'b11001110;
DRAM[36981] = 8'b11011110;
DRAM[36982] = 8'b11101000;
DRAM[36983] = 8'b11101001;
DRAM[36984] = 8'b11100100;
DRAM[36985] = 8'b11100010;
DRAM[36986] = 8'b11011111;
DRAM[36987] = 8'b11011110;
DRAM[36988] = 8'b11100000;
DRAM[36989] = 8'b11100011;
DRAM[36990] = 8'b11100011;
DRAM[36991] = 8'b11100011;
DRAM[36992] = 8'b11100111;
DRAM[36993] = 8'b11100110;
DRAM[36994] = 8'b11100011;
DRAM[36995] = 8'b11011001;
DRAM[36996] = 8'b11011000;
DRAM[36997] = 8'b11101100;
DRAM[36998] = 8'b11110100;
DRAM[36999] = 8'b11100110;
DRAM[37000] = 8'b11101011;
DRAM[37001] = 8'b11100011;
DRAM[37002] = 8'b11010111;
DRAM[37003] = 8'b11001100;
DRAM[37004] = 8'b11000101;
DRAM[37005] = 8'b11000000;
DRAM[37006] = 8'b10111011;
DRAM[37007] = 8'b10111000;
DRAM[37008] = 8'b10100000;
DRAM[37009] = 8'b10011101;
DRAM[37010] = 8'b10011000;
DRAM[37011] = 8'b10010110;
DRAM[37012] = 8'b10010111;
DRAM[37013] = 8'b10011011;
DRAM[37014] = 8'b10100001;
DRAM[37015] = 8'b10100110;
DRAM[37016] = 8'b10101100;
DRAM[37017] = 8'b10110100;
DRAM[37018] = 8'b10111111;
DRAM[37019] = 8'b10110101;
DRAM[37020] = 8'b10101110;
DRAM[37021] = 8'b11001111;
DRAM[37022] = 8'b11101001;
DRAM[37023] = 8'b11011101;
DRAM[37024] = 8'b11000011;
DRAM[37025] = 8'b11001011;
DRAM[37026] = 8'b11010110;
DRAM[37027] = 8'b11100000;
DRAM[37028] = 8'b11101010;
DRAM[37029] = 8'b11110010;
DRAM[37030] = 8'b11110100;
DRAM[37031] = 8'b11110011;
DRAM[37032] = 8'b11110011;
DRAM[37033] = 8'b11101111;
DRAM[37034] = 8'b11101000;
DRAM[37035] = 8'b11100111;
DRAM[37036] = 8'b11101101;
DRAM[37037] = 8'b11101100;
DRAM[37038] = 8'b11010101;
DRAM[37039] = 8'b10111010;
DRAM[37040] = 8'b10100110;
DRAM[37041] = 8'b10101010;
DRAM[37042] = 8'b10110010;
DRAM[37043] = 8'b10111101;
DRAM[37044] = 8'b11001000;
DRAM[37045] = 8'b11001011;
DRAM[37046] = 8'b11000100;
DRAM[37047] = 8'b10111010;
DRAM[37048] = 8'b10110110;
DRAM[37049] = 8'b10111001;
DRAM[37050] = 8'b10111010;
DRAM[37051] = 8'b10111010;
DRAM[37052] = 8'b10111100;
DRAM[37053] = 8'b10111011;
DRAM[37054] = 8'b10101111;
DRAM[37055] = 8'b10100001;
DRAM[37056] = 8'b10100010;
DRAM[37057] = 8'b10011010;
DRAM[37058] = 8'b10010111;
DRAM[37059] = 8'b10011101;
DRAM[37060] = 8'b10100110;
DRAM[37061] = 8'b10101101;
DRAM[37062] = 8'b10110100;
DRAM[37063] = 8'b10111010;
DRAM[37064] = 8'b11011100;
DRAM[37065] = 8'b11011100;
DRAM[37066] = 8'b11100000;
DRAM[37067] = 8'b11011010;
DRAM[37068] = 8'b11001110;
DRAM[37069] = 8'b11001011;
DRAM[37070] = 8'b11000010;
DRAM[37071] = 8'b10101110;
DRAM[37072] = 8'b10100010;
DRAM[37073] = 8'b10011010;
DRAM[37074] = 8'b10010011;
DRAM[37075] = 8'b10010001;
DRAM[37076] = 8'b10001111;
DRAM[37077] = 8'b10001100;
DRAM[37078] = 8'b10001100;
DRAM[37079] = 8'b10001111;
DRAM[37080] = 8'b10001110;
DRAM[37081] = 8'b10001101;
DRAM[37082] = 8'b10001100;
DRAM[37083] = 8'b10001011;
DRAM[37084] = 8'b10001011;
DRAM[37085] = 8'b10001011;
DRAM[37086] = 8'b10001011;
DRAM[37087] = 8'b10001100;
DRAM[37088] = 8'b10001000;
DRAM[37089] = 8'b10001000;
DRAM[37090] = 8'b10001000;
DRAM[37091] = 8'b10001000;
DRAM[37092] = 8'b10001000;
DRAM[37093] = 8'b10000110;
DRAM[37094] = 8'b10000101;
DRAM[37095] = 8'b10000101;
DRAM[37096] = 8'b10000110;
DRAM[37097] = 8'b10000110;
DRAM[37098] = 8'b10000100;
DRAM[37099] = 8'b10000011;
DRAM[37100] = 8'b10000010;
DRAM[37101] = 8'b10000001;
DRAM[37102] = 8'b10000001;
DRAM[37103] = 8'b10000010;
DRAM[37104] = 8'b10000001;
DRAM[37105] = 8'b10000000;
DRAM[37106] = 8'b1111110;
DRAM[37107] = 8'b1111100;
DRAM[37108] = 8'b1111011;
DRAM[37109] = 8'b1111011;
DRAM[37110] = 8'b1111100;
DRAM[37111] = 8'b1111100;
DRAM[37112] = 8'b1111011;
DRAM[37113] = 8'b1111011;
DRAM[37114] = 8'b1111011;
DRAM[37115] = 8'b1111011;
DRAM[37116] = 8'b1111011;
DRAM[37117] = 8'b1111011;
DRAM[37118] = 8'b1111011;
DRAM[37119] = 8'b1111011;
DRAM[37120] = 8'b10011000;
DRAM[37121] = 8'b10011000;
DRAM[37122] = 8'b10011001;
DRAM[37123] = 8'b10011010;
DRAM[37124] = 8'b10011011;
DRAM[37125] = 8'b10011011;
DRAM[37126] = 8'b10011100;
DRAM[37127] = 8'b10011100;
DRAM[37128] = 8'b10011101;
DRAM[37129] = 8'b10011101;
DRAM[37130] = 8'b10011110;
DRAM[37131] = 8'b10011110;
DRAM[37132] = 8'b10011110;
DRAM[37133] = 8'b10011110;
DRAM[37134] = 8'b10011111;
DRAM[37135] = 8'b10011111;
DRAM[37136] = 8'b10100000;
DRAM[37137] = 8'b10100000;
DRAM[37138] = 8'b10011111;
DRAM[37139] = 8'b10011111;
DRAM[37140] = 8'b10100000;
DRAM[37141] = 8'b10100000;
DRAM[37142] = 8'b10100001;
DRAM[37143] = 8'b10100010;
DRAM[37144] = 8'b10100000;
DRAM[37145] = 8'b10100000;
DRAM[37146] = 8'b10100000;
DRAM[37147] = 8'b10100000;
DRAM[37148] = 8'b10100001;
DRAM[37149] = 8'b10100010;
DRAM[37150] = 8'b10100011;
DRAM[37151] = 8'b10100100;
DRAM[37152] = 8'b10100100;
DRAM[37153] = 8'b10100101;
DRAM[37154] = 8'b10100110;
DRAM[37155] = 8'b10100111;
DRAM[37156] = 8'b10101000;
DRAM[37157] = 8'b10100111;
DRAM[37158] = 8'b10100111;
DRAM[37159] = 8'b10100111;
DRAM[37160] = 8'b10100101;
DRAM[37161] = 8'b10100100;
DRAM[37162] = 8'b10100100;
DRAM[37163] = 8'b10100011;
DRAM[37164] = 8'b10100011;
DRAM[37165] = 8'b10100100;
DRAM[37166] = 8'b10100100;
DRAM[37167] = 8'b10100101;
DRAM[37168] = 8'b10100001;
DRAM[37169] = 8'b10100110;
DRAM[37170] = 8'b10101010;
DRAM[37171] = 8'b10101011;
DRAM[37172] = 8'b10101010;
DRAM[37173] = 8'b10101110;
DRAM[37174] = 8'b10110110;
DRAM[37175] = 8'b10111110;
DRAM[37176] = 8'b11011001;
DRAM[37177] = 8'b11100110;
DRAM[37178] = 8'b11110100;
DRAM[37179] = 8'b11111011;
DRAM[37180] = 8'b11111101;
DRAM[37181] = 8'b11111100;
DRAM[37182] = 8'b11110111;
DRAM[37183] = 8'b11110000;
DRAM[37184] = 8'b11011110;
DRAM[37185] = 8'b11010101;
DRAM[37186] = 8'b11001000;
DRAM[37187] = 8'b10111110;
DRAM[37188] = 8'b10111000;
DRAM[37189] = 8'b10110100;
DRAM[37190] = 8'b10110000;
DRAM[37191] = 8'b10101100;
DRAM[37192] = 8'b10101001;
DRAM[37193] = 8'b10100111;
DRAM[37194] = 8'b10100101;
DRAM[37195] = 8'b10100100;
DRAM[37196] = 8'b10100100;
DRAM[37197] = 8'b10100000;
DRAM[37198] = 8'b10011001;
DRAM[37199] = 8'b10010100;
DRAM[37200] = 8'b10100010;
DRAM[37201] = 8'b10100010;
DRAM[37202] = 8'b10100000;
DRAM[37203] = 8'b10100100;
DRAM[37204] = 8'b10101101;
DRAM[37205] = 8'b10101011;
DRAM[37206] = 8'b10101001;
DRAM[37207] = 8'b10110001;
DRAM[37208] = 8'b10101000;
DRAM[37209] = 8'b10110000;
DRAM[37210] = 8'b10111001;
DRAM[37211] = 8'b10111110;
DRAM[37212] = 8'b10111110;
DRAM[37213] = 8'b10111011;
DRAM[37214] = 8'b10111010;
DRAM[37215] = 8'b10111011;
DRAM[37216] = 8'b10110100;
DRAM[37217] = 8'b10111011;
DRAM[37218] = 8'b11000001;
DRAM[37219] = 8'b11000001;
DRAM[37220] = 8'b10111011;
DRAM[37221] = 8'b10110111;
DRAM[37222] = 8'b10111000;
DRAM[37223] = 8'b10111100;
DRAM[37224] = 8'b10101001;
DRAM[37225] = 8'b10110011;
DRAM[37226] = 8'b10111001;
DRAM[37227] = 8'b10110111;
DRAM[37228] = 8'b10110100;
DRAM[37229] = 8'b10110111;
DRAM[37230] = 8'b10111011;
DRAM[37231] = 8'b10111100;
DRAM[37232] = 8'b10100011;
DRAM[37233] = 8'b10110110;
DRAM[37234] = 8'b11000101;
DRAM[37235] = 8'b11001000;
DRAM[37236] = 8'b11001101;
DRAM[37237] = 8'b11011010;
DRAM[37238] = 8'b11100011;
DRAM[37239] = 8'b11100011;
DRAM[37240] = 8'b11100110;
DRAM[37241] = 8'b11100101;
DRAM[37242] = 8'b11100010;
DRAM[37243] = 8'b11011110;
DRAM[37244] = 8'b11011011;
DRAM[37245] = 8'b11011011;
DRAM[37246] = 8'b11011101;
DRAM[37247] = 8'b11011111;
DRAM[37248] = 8'b11101001;
DRAM[37249] = 8'b11011010;
DRAM[37250] = 8'b11010011;
DRAM[37251] = 8'b11010100;
DRAM[37252] = 8'b11010110;
DRAM[37253] = 8'b11011111;
DRAM[37254] = 8'b11100011;
DRAM[37255] = 8'b11011000;
DRAM[37256] = 8'b11010010;
DRAM[37257] = 8'b11000110;
DRAM[37258] = 8'b10110101;
DRAM[37259] = 8'b10100111;
DRAM[37260] = 8'b10011111;
DRAM[37261] = 8'b10011010;
DRAM[37262] = 8'b10010110;
DRAM[37263] = 8'b10010011;
DRAM[37264] = 8'b10001011;
DRAM[37265] = 8'b10001000;
DRAM[37266] = 8'b10000011;
DRAM[37267] = 8'b10000000;
DRAM[37268] = 8'b10000000;
DRAM[37269] = 8'b10000100;
DRAM[37270] = 8'b10001001;
DRAM[37271] = 8'b10001101;
DRAM[37272] = 8'b10001110;
DRAM[37273] = 8'b10010001;
DRAM[37274] = 8'b10011000;
DRAM[37275] = 8'b10011101;
DRAM[37276] = 8'b10101000;
DRAM[37277] = 8'b10111111;
DRAM[37278] = 8'b11000110;
DRAM[37279] = 8'b10111001;
DRAM[37280] = 8'b10111100;
DRAM[37281] = 8'b11000111;
DRAM[37282] = 8'b11010100;
DRAM[37283] = 8'b11011111;
DRAM[37284] = 8'b11101001;
DRAM[37285] = 8'b11110001;
DRAM[37286] = 8'b11110011;
DRAM[37287] = 8'b11110010;
DRAM[37288] = 8'b11110101;
DRAM[37289] = 8'b11110011;
DRAM[37290] = 8'b11101101;
DRAM[37291] = 8'b11101100;
DRAM[37292] = 8'b11110100;
DRAM[37293] = 8'b11110101;
DRAM[37294] = 8'b11100010;
DRAM[37295] = 8'b11001010;
DRAM[37296] = 8'b10100101;
DRAM[37297] = 8'b10101000;
DRAM[37298] = 8'b10101100;
DRAM[37299] = 8'b10110011;
DRAM[37300] = 8'b10111100;
DRAM[37301] = 8'b11000011;
DRAM[37302] = 8'b11000110;
DRAM[37303] = 8'b11000110;
DRAM[37304] = 8'b10111100;
DRAM[37305] = 8'b10111101;
DRAM[37306] = 8'b10111010;
DRAM[37307] = 8'b10111000;
DRAM[37308] = 8'b10111010;
DRAM[37309] = 8'b10111011;
DRAM[37310] = 8'b10110010;
DRAM[37311] = 8'b10100111;
DRAM[37312] = 8'b10011010;
DRAM[37313] = 8'b10010110;
DRAM[37314] = 8'b10010111;
DRAM[37315] = 8'b10100000;
DRAM[37316] = 8'b10101101;
DRAM[37317] = 8'b10111011;
DRAM[37318] = 8'b11001001;
DRAM[37319] = 8'b11010100;
DRAM[37320] = 8'b11011111;
DRAM[37321] = 8'b11100001;
DRAM[37322] = 8'b11100111;
DRAM[37323] = 8'b11100001;
DRAM[37324] = 8'b11010001;
DRAM[37325] = 8'b11000111;
DRAM[37326] = 8'b10110110;
DRAM[37327] = 8'b10011100;
DRAM[37328] = 8'b10100100;
DRAM[37329] = 8'b10011100;
DRAM[37330] = 8'b10010101;
DRAM[37331] = 8'b10010011;
DRAM[37332] = 8'b10010001;
DRAM[37333] = 8'b10001101;
DRAM[37334] = 8'b10001100;
DRAM[37335] = 8'b10001110;
DRAM[37336] = 8'b10001110;
DRAM[37337] = 8'b10001101;
DRAM[37338] = 8'b10001100;
DRAM[37339] = 8'b10001100;
DRAM[37340] = 8'b10001011;
DRAM[37341] = 8'b10001011;
DRAM[37342] = 8'b10001100;
DRAM[37343] = 8'b10001100;
DRAM[37344] = 8'b10001001;
DRAM[37345] = 8'b10001001;
DRAM[37346] = 8'b10001001;
DRAM[37347] = 8'b10001000;
DRAM[37348] = 8'b10000111;
DRAM[37349] = 8'b10000110;
DRAM[37350] = 8'b10000101;
DRAM[37351] = 8'b10000100;
DRAM[37352] = 8'b10000101;
DRAM[37353] = 8'b10000101;
DRAM[37354] = 8'b10000011;
DRAM[37355] = 8'b10000010;
DRAM[37356] = 8'b10000001;
DRAM[37357] = 8'b10000001;
DRAM[37358] = 8'b10000001;
DRAM[37359] = 8'b10000001;
DRAM[37360] = 8'b10000001;
DRAM[37361] = 8'b10000000;
DRAM[37362] = 8'b1111110;
DRAM[37363] = 8'b1111100;
DRAM[37364] = 8'b1111011;
DRAM[37365] = 8'b1111011;
DRAM[37366] = 8'b1111100;
DRAM[37367] = 8'b1111100;
DRAM[37368] = 8'b1111011;
DRAM[37369] = 8'b1111011;
DRAM[37370] = 8'b1111011;
DRAM[37371] = 8'b1111011;
DRAM[37372] = 8'b1111011;
DRAM[37373] = 8'b1111011;
DRAM[37374] = 8'b1111011;
DRAM[37375] = 8'b1111011;
DRAM[37376] = 8'b10011000;
DRAM[37377] = 8'b10011001;
DRAM[37378] = 8'b10011001;
DRAM[37379] = 8'b10011010;
DRAM[37380] = 8'b10011011;
DRAM[37381] = 8'b10011100;
DRAM[37382] = 8'b10011100;
DRAM[37383] = 8'b10011100;
DRAM[37384] = 8'b10011101;
DRAM[37385] = 8'b10011101;
DRAM[37386] = 8'b10011101;
DRAM[37387] = 8'b10011110;
DRAM[37388] = 8'b10011110;
DRAM[37389] = 8'b10011111;
DRAM[37390] = 8'b10011111;
DRAM[37391] = 8'b10011111;
DRAM[37392] = 8'b10100000;
DRAM[37393] = 8'b10100000;
DRAM[37394] = 8'b10011111;
DRAM[37395] = 8'b10011111;
DRAM[37396] = 8'b10100000;
DRAM[37397] = 8'b10100001;
DRAM[37398] = 8'b10100010;
DRAM[37399] = 8'b10100010;
DRAM[37400] = 8'b10100010;
DRAM[37401] = 8'b10100010;
DRAM[37402] = 8'b10100001;
DRAM[37403] = 8'b10100001;
DRAM[37404] = 8'b10100001;
DRAM[37405] = 8'b10100010;
DRAM[37406] = 8'b10100010;
DRAM[37407] = 8'b10100011;
DRAM[37408] = 8'b10100100;
DRAM[37409] = 8'b10100100;
DRAM[37410] = 8'b10100101;
DRAM[37411] = 8'b10100110;
DRAM[37412] = 8'b10100111;
DRAM[37413] = 8'b10100110;
DRAM[37414] = 8'b10100110;
DRAM[37415] = 8'b10100110;
DRAM[37416] = 8'b10100101;
DRAM[37417] = 8'b10100100;
DRAM[37418] = 8'b10100100;
DRAM[37419] = 8'b10100011;
DRAM[37420] = 8'b10100011;
DRAM[37421] = 8'b10100100;
DRAM[37422] = 8'b10100100;
DRAM[37423] = 8'b10100101;
DRAM[37424] = 8'b10101000;
DRAM[37425] = 8'b10101000;
DRAM[37426] = 8'b10100101;
DRAM[37427] = 8'b10100010;
DRAM[37428] = 8'b10100111;
DRAM[37429] = 8'b10111000;
DRAM[37430] = 8'b11010010;
DRAM[37431] = 8'b11100110;
DRAM[37432] = 8'b11110101;
DRAM[37433] = 8'b11111010;
DRAM[37434] = 8'b11111100;
DRAM[37435] = 8'b11111100;
DRAM[37436] = 8'b11111100;
DRAM[37437] = 8'b11111011;
DRAM[37438] = 8'b11110101;
DRAM[37439] = 8'b11101110;
DRAM[37440] = 8'b11011110;
DRAM[37441] = 8'b11010101;
DRAM[37442] = 8'b11001000;
DRAM[37443] = 8'b10111110;
DRAM[37444] = 8'b10111001;
DRAM[37445] = 8'b10110110;
DRAM[37446] = 8'b10110010;
DRAM[37447] = 8'b10110000;
DRAM[37448] = 8'b10101010;
DRAM[37449] = 8'b10101010;
DRAM[37450] = 8'b10101001;
DRAM[37451] = 8'b10101001;
DRAM[37452] = 8'b10100111;
DRAM[37453] = 8'b10100110;
DRAM[37454] = 8'b10100100;
DRAM[37455] = 8'b10100010;
DRAM[37456] = 8'b10110010;
DRAM[37457] = 8'b10100100;
DRAM[37458] = 8'b10100010;
DRAM[37459] = 8'b10101000;
DRAM[37460] = 8'b10101001;
DRAM[37461] = 8'b10101000;
DRAM[37462] = 8'b10100011;
DRAM[37463] = 8'b10011000;
DRAM[37464] = 8'b10100010;
DRAM[37465] = 8'b10101000;
DRAM[37466] = 8'b10101110;
DRAM[37467] = 8'b10110001;
DRAM[37468] = 8'b10110010;
DRAM[37469] = 8'b10110110;
DRAM[37470] = 8'b10111110;
DRAM[37471] = 8'b11000101;
DRAM[37472] = 8'b10111111;
DRAM[37473] = 8'b10111010;
DRAM[37474] = 8'b10111000;
DRAM[37475] = 8'b10111100;
DRAM[37476] = 8'b11000001;
DRAM[37477] = 8'b11000000;
DRAM[37478] = 8'b10110101;
DRAM[37479] = 8'b10101011;
DRAM[37480] = 8'b10110101;
DRAM[37481] = 8'b11000000;
DRAM[37482] = 8'b11000000;
DRAM[37483] = 8'b10110101;
DRAM[37484] = 8'b10110101;
DRAM[37485] = 8'b10111101;
DRAM[37486] = 8'b10110111;
DRAM[37487] = 8'b10100110;
DRAM[37488] = 8'b10101100;
DRAM[37489] = 8'b10111111;
DRAM[37490] = 8'b11001111;
DRAM[37491] = 8'b11010001;
DRAM[37492] = 8'b11010000;
DRAM[37493] = 8'b11010101;
DRAM[37494] = 8'b11011010;
DRAM[37495] = 8'b11011010;
DRAM[37496] = 8'b11100000;
DRAM[37497] = 8'b11100010;
DRAM[37498] = 8'b11100001;
DRAM[37499] = 8'b11011011;
DRAM[37500] = 8'b11010011;
DRAM[37501] = 8'b11010010;
DRAM[37502] = 8'b11011000;
DRAM[37503] = 8'b11011111;
DRAM[37504] = 8'b11011101;
DRAM[37505] = 8'b11000100;
DRAM[37506] = 8'b10111101;
DRAM[37507] = 8'b11001000;
DRAM[37508] = 8'b11001110;
DRAM[37509] = 8'b11010011;
DRAM[37510] = 8'b11010010;
DRAM[37511] = 8'b11001011;
DRAM[37512] = 8'b10110100;
DRAM[37513] = 8'b10100100;
DRAM[37514] = 8'b10001111;
DRAM[37515] = 8'b1111110;
DRAM[37516] = 8'b1110110;
DRAM[37517] = 8'b1110100;
DRAM[37518] = 8'b1110010;
DRAM[37519] = 8'b1110001;
DRAM[37520] = 8'b1110101;
DRAM[37521] = 8'b1110011;
DRAM[37522] = 8'b1101111;
DRAM[37523] = 8'b1101101;
DRAM[37524] = 8'b1101110;
DRAM[37525] = 8'b1110010;
DRAM[37526] = 8'b1110110;
DRAM[37527] = 8'b1111010;
DRAM[37528] = 8'b1111000;
DRAM[37529] = 8'b1111001;
DRAM[37530] = 8'b1111001;
DRAM[37531] = 8'b10000010;
DRAM[37532] = 8'b10010101;
DRAM[37533] = 8'b10011110;
DRAM[37534] = 8'b10100100;
DRAM[37535] = 8'b10101110;
DRAM[37536] = 8'b11000011;
DRAM[37537] = 8'b11010000;
DRAM[37538] = 8'b11011110;
DRAM[37539] = 8'b11100100;
DRAM[37540] = 8'b11101001;
DRAM[37541] = 8'b11101110;
DRAM[37542] = 8'b11110000;
DRAM[37543] = 8'b11101111;
DRAM[37544] = 8'b11110111;
DRAM[37545] = 8'b11110111;
DRAM[37546] = 8'b11110011;
DRAM[37547] = 8'b11110001;
DRAM[37548] = 8'b11110111;
DRAM[37549] = 8'b11111010;
DRAM[37550] = 8'b11101100;
DRAM[37551] = 8'b11011000;
DRAM[37552] = 8'b10111111;
DRAM[37553] = 8'b10111101;
DRAM[37554] = 8'b10111011;
DRAM[37555] = 8'b10111000;
DRAM[37556] = 8'b10110101;
DRAM[37557] = 8'b10110100;
DRAM[37558] = 8'b10110101;
DRAM[37559] = 8'b10111000;
DRAM[37560] = 8'b11000001;
DRAM[37561] = 8'b10111110;
DRAM[37562] = 8'b10111000;
DRAM[37563] = 8'b10110101;
DRAM[37564] = 8'b10110111;
DRAM[37565] = 8'b10111010;
DRAM[37566] = 8'b10110101;
DRAM[37567] = 8'b10101110;
DRAM[37568] = 8'b10011110;
DRAM[37569] = 8'b10011011;
DRAM[37570] = 8'b10011011;
DRAM[37571] = 8'b10100011;
DRAM[37572] = 8'b10101101;
DRAM[37573] = 8'b10111011;
DRAM[37574] = 8'b11001101;
DRAM[37575] = 8'b11011100;
DRAM[37576] = 8'b11100110;
DRAM[37577] = 8'b11100010;
DRAM[37578] = 8'b11011110;
DRAM[37579] = 8'b11010001;
DRAM[37580] = 8'b11000001;
DRAM[37581] = 8'b10111100;
DRAM[37582] = 8'b10110100;
DRAM[37583] = 8'b10100001;
DRAM[37584] = 8'b10100010;
DRAM[37585] = 8'b10011010;
DRAM[37586] = 8'b10010100;
DRAM[37587] = 8'b10010011;
DRAM[37588] = 8'b10010001;
DRAM[37589] = 8'b10001110;
DRAM[37590] = 8'b10001101;
DRAM[37591] = 8'b10001111;
DRAM[37592] = 8'b10001110;
DRAM[37593] = 8'b10001110;
DRAM[37594] = 8'b10001101;
DRAM[37595] = 8'b10001100;
DRAM[37596] = 8'b10001011;
DRAM[37597] = 8'b10001011;
DRAM[37598] = 8'b10001100;
DRAM[37599] = 8'b10001100;
DRAM[37600] = 8'b10001010;
DRAM[37601] = 8'b10001010;
DRAM[37602] = 8'b10001001;
DRAM[37603] = 8'b10001001;
DRAM[37604] = 8'b10000111;
DRAM[37605] = 8'b10000101;
DRAM[37606] = 8'b10000011;
DRAM[37607] = 8'b10000010;
DRAM[37608] = 8'b10000100;
DRAM[37609] = 8'b10000011;
DRAM[37610] = 8'b10000010;
DRAM[37611] = 8'b10000001;
DRAM[37612] = 8'b10000000;
DRAM[37613] = 8'b10000000;
DRAM[37614] = 8'b10000000;
DRAM[37615] = 8'b10000000;
DRAM[37616] = 8'b10000000;
DRAM[37617] = 8'b1111111;
DRAM[37618] = 8'b1111101;
DRAM[37619] = 8'b1111100;
DRAM[37620] = 8'b1111011;
DRAM[37621] = 8'b1111011;
DRAM[37622] = 8'b1111100;
DRAM[37623] = 8'b1111101;
DRAM[37624] = 8'b1111011;
DRAM[37625] = 8'b1111011;
DRAM[37626] = 8'b1111011;
DRAM[37627] = 8'b1111011;
DRAM[37628] = 8'b1111011;
DRAM[37629] = 8'b1111011;
DRAM[37630] = 8'b1111011;
DRAM[37631] = 8'b1111011;
DRAM[37632] = 8'b10011001;
DRAM[37633] = 8'b10011001;
DRAM[37634] = 8'b10011010;
DRAM[37635] = 8'b10011010;
DRAM[37636] = 8'b10011011;
DRAM[37637] = 8'b10011100;
DRAM[37638] = 8'b10011101;
DRAM[37639] = 8'b10011101;
DRAM[37640] = 8'b10011100;
DRAM[37641] = 8'b10011100;
DRAM[37642] = 8'b10011101;
DRAM[37643] = 8'b10011110;
DRAM[37644] = 8'b10011110;
DRAM[37645] = 8'b10011111;
DRAM[37646] = 8'b10100000;
DRAM[37647] = 8'b10100000;
DRAM[37648] = 8'b10100001;
DRAM[37649] = 8'b10100000;
DRAM[37650] = 8'b10100000;
DRAM[37651] = 8'b10100000;
DRAM[37652] = 8'b10100000;
DRAM[37653] = 8'b10100001;
DRAM[37654] = 8'b10100010;
DRAM[37655] = 8'b10100011;
DRAM[37656] = 8'b10100100;
DRAM[37657] = 8'b10100011;
DRAM[37658] = 8'b10100011;
DRAM[37659] = 8'b10100010;
DRAM[37660] = 8'b10100010;
DRAM[37661] = 8'b10100010;
DRAM[37662] = 8'b10100010;
DRAM[37663] = 8'b10100011;
DRAM[37664] = 8'b10100100;
DRAM[37665] = 8'b10100100;
DRAM[37666] = 8'b10100101;
DRAM[37667] = 8'b10100110;
DRAM[37668] = 8'b10100110;
DRAM[37669] = 8'b10100101;
DRAM[37670] = 8'b10100101;
DRAM[37671] = 8'b10100100;
DRAM[37672] = 8'b10100101;
DRAM[37673] = 8'b10100100;
DRAM[37674] = 8'b10100100;
DRAM[37675] = 8'b10100011;
DRAM[37676] = 8'b10100011;
DRAM[37677] = 8'b10100100;
DRAM[37678] = 8'b10100100;
DRAM[37679] = 8'b10100101;
DRAM[37680] = 8'b10101011;
DRAM[37681] = 8'b10101000;
DRAM[37682] = 8'b10100100;
DRAM[37683] = 8'b10100010;
DRAM[37684] = 8'b10101011;
DRAM[37685] = 8'b11000100;
DRAM[37686] = 8'b11100110;
DRAM[37687] = 8'b11111110;
DRAM[37688] = 8'b11111100;
DRAM[37689] = 8'b11111100;
DRAM[37690] = 8'b11111010;
DRAM[37691] = 8'b11111000;
DRAM[37692] = 8'b11111010;
DRAM[37693] = 8'b11111011;
DRAM[37694] = 8'b11110101;
DRAM[37695] = 8'b11101011;
DRAM[37696] = 8'b11011101;
DRAM[37697] = 8'b11010101;
DRAM[37698] = 8'b11001011;
DRAM[37699] = 8'b11000010;
DRAM[37700] = 8'b10111110;
DRAM[37701] = 8'b10111010;
DRAM[37702] = 8'b10110101;
DRAM[37703] = 8'b10110010;
DRAM[37704] = 8'b10101110;
DRAM[37705] = 8'b10101111;
DRAM[37706] = 8'b10101111;
DRAM[37707] = 8'b10101101;
DRAM[37708] = 8'b10101011;
DRAM[37709] = 8'b10101010;
DRAM[37710] = 8'b10101011;
DRAM[37711] = 8'b10101100;
DRAM[37712] = 8'b10101001;
DRAM[37713] = 8'b10100001;
DRAM[37714] = 8'b10101100;
DRAM[37715] = 8'b10110010;
DRAM[37716] = 8'b10100110;
DRAM[37717] = 8'b10101001;
DRAM[37718] = 8'b10110011;
DRAM[37719] = 8'b10101100;
DRAM[37720] = 8'b10100111;
DRAM[37721] = 8'b10101001;
DRAM[37722] = 8'b10101001;
DRAM[37723] = 8'b10100111;
DRAM[37724] = 8'b10101000;
DRAM[37725] = 8'b10101110;
DRAM[37726] = 8'b10111010;
DRAM[37727] = 8'b11000100;
DRAM[37728] = 8'b11001000;
DRAM[37729] = 8'b10111100;
DRAM[37730] = 8'b10110000;
DRAM[37731] = 8'b10110001;
DRAM[37732] = 8'b10111010;
DRAM[37733] = 8'b11000000;
DRAM[37734] = 8'b10111011;
DRAM[37735] = 8'b10110100;
DRAM[37736] = 8'b11000101;
DRAM[37737] = 8'b10111100;
DRAM[37738] = 8'b10111100;
DRAM[37739] = 8'b11000110;
DRAM[37740] = 8'b11000110;
DRAM[37741] = 8'b10111000;
DRAM[37742] = 8'b10101011;
DRAM[37743] = 8'b10101000;
DRAM[37744] = 8'b10111010;
DRAM[37745] = 8'b11001001;
DRAM[37746] = 8'b11010101;
DRAM[37747] = 8'b11010011;
DRAM[37748] = 8'b11001111;
DRAM[37749] = 8'b11010001;
DRAM[37750] = 8'b11010111;
DRAM[37751] = 8'b11011010;
DRAM[37752] = 8'b11011110;
DRAM[37753] = 8'b11100010;
DRAM[37754] = 8'b11100010;
DRAM[37755] = 8'b11011010;
DRAM[37756] = 8'b11001110;
DRAM[37757] = 8'b11001010;
DRAM[37758] = 8'b11010001;
DRAM[37759] = 8'b11011001;
DRAM[37760] = 8'b11010011;
DRAM[37761] = 8'b10111110;
DRAM[37762] = 8'b10110100;
DRAM[37763] = 8'b10111000;
DRAM[37764] = 8'b10111001;
DRAM[37765] = 8'b10111101;
DRAM[37766] = 8'b10111010;
DRAM[37767] = 8'b10101101;
DRAM[37768] = 8'b10011010;
DRAM[37769] = 8'b10001011;
DRAM[37770] = 8'b1110110;
DRAM[37771] = 8'b1100111;
DRAM[37772] = 8'b1100010;
DRAM[37773] = 8'b1100100;
DRAM[37774] = 8'b1100110;
DRAM[37775] = 8'b1101000;
DRAM[37776] = 8'b1101011;
DRAM[37777] = 8'b1101001;
DRAM[37778] = 8'b1100111;
DRAM[37779] = 8'b1100110;
DRAM[37780] = 8'b1101000;
DRAM[37781] = 8'b1101100;
DRAM[37782] = 8'b1110001;
DRAM[37783] = 8'b1110011;
DRAM[37784] = 8'b1110011;
DRAM[37785] = 8'b1111010;
DRAM[37786] = 8'b1110101;
DRAM[37787] = 8'b1110101;
DRAM[37788] = 8'b1111010;
DRAM[37789] = 8'b1110111;
DRAM[37790] = 8'b10001010;
DRAM[37791] = 8'b10110111;
DRAM[37792] = 8'b11000010;
DRAM[37793] = 8'b11010010;
DRAM[37794] = 8'b11011111;
DRAM[37795] = 8'b11100000;
DRAM[37796] = 8'b11100001;
DRAM[37797] = 8'b11101000;
DRAM[37798] = 8'b11101110;
DRAM[37799] = 8'b11101111;
DRAM[37800] = 8'b11110101;
DRAM[37801] = 8'b11111000;
DRAM[37802] = 8'b11110101;
DRAM[37803] = 8'b11110000;
DRAM[37804] = 8'b11110011;
DRAM[37805] = 8'b11110110;
DRAM[37806] = 8'b11101100;
DRAM[37807] = 8'b11011110;
DRAM[37808] = 8'b10111011;
DRAM[37809] = 8'b10110111;
DRAM[37810] = 8'b10110111;
DRAM[37811] = 8'b10111010;
DRAM[37812] = 8'b10111101;
DRAM[37813] = 8'b10111101;
DRAM[37814] = 8'b10111100;
DRAM[37815] = 8'b10111101;
DRAM[37816] = 8'b10111101;
DRAM[37817] = 8'b10111001;
DRAM[37818] = 8'b10110011;
DRAM[37819] = 8'b10110010;
DRAM[37820] = 8'b10110110;
DRAM[37821] = 8'b10111001;
DRAM[37822] = 8'b10110110;
DRAM[37823] = 8'b10110001;
DRAM[37824] = 8'b10100110;
DRAM[37825] = 8'b10100011;
DRAM[37826] = 8'b10100011;
DRAM[37827] = 8'b10100111;
DRAM[37828] = 8'b10101110;
DRAM[37829] = 8'b10111011;
DRAM[37830] = 8'b11001110;
DRAM[37831] = 8'b11011111;
DRAM[37832] = 8'b11101000;
DRAM[37833] = 8'b11100010;
DRAM[37834] = 8'b11011100;
DRAM[37835] = 8'b11001101;
DRAM[37836] = 8'b10111101;
DRAM[37837] = 8'b10111011;
DRAM[37838] = 8'b10110111;
DRAM[37839] = 8'b10100110;
DRAM[37840] = 8'b10011101;
DRAM[37841] = 8'b10010111;
DRAM[37842] = 8'b10010010;
DRAM[37843] = 8'b10010010;
DRAM[37844] = 8'b10010001;
DRAM[37845] = 8'b10001111;
DRAM[37846] = 8'b10001110;
DRAM[37847] = 8'b10010001;
DRAM[37848] = 8'b10001111;
DRAM[37849] = 8'b10001110;
DRAM[37850] = 8'b10001101;
DRAM[37851] = 8'b10001100;
DRAM[37852] = 8'b10001100;
DRAM[37853] = 8'b10001100;
DRAM[37854] = 8'b10001100;
DRAM[37855] = 8'b10001101;
DRAM[37856] = 8'b10001011;
DRAM[37857] = 8'b10001011;
DRAM[37858] = 8'b10001010;
DRAM[37859] = 8'b10001001;
DRAM[37860] = 8'b10000111;
DRAM[37861] = 8'b10000101;
DRAM[37862] = 8'b10000011;
DRAM[37863] = 8'b10000001;
DRAM[37864] = 8'b10000010;
DRAM[37865] = 8'b10000010;
DRAM[37866] = 8'b10000000;
DRAM[37867] = 8'b10000000;
DRAM[37868] = 8'b1111111;
DRAM[37869] = 8'b1111111;
DRAM[37870] = 8'b1111111;
DRAM[37871] = 8'b10000000;
DRAM[37872] = 8'b10000000;
DRAM[37873] = 8'b1111111;
DRAM[37874] = 8'b1111101;
DRAM[37875] = 8'b1111100;
DRAM[37876] = 8'b1111011;
DRAM[37877] = 8'b1111100;
DRAM[37878] = 8'b1111101;
DRAM[37879] = 8'b1111101;
DRAM[37880] = 8'b1111100;
DRAM[37881] = 8'b1111100;
DRAM[37882] = 8'b1111100;
DRAM[37883] = 8'b1111100;
DRAM[37884] = 8'b1111100;
DRAM[37885] = 8'b1111100;
DRAM[37886] = 8'b1111100;
DRAM[37887] = 8'b1111100;
DRAM[37888] = 8'b10011001;
DRAM[37889] = 8'b10011001;
DRAM[37890] = 8'b10011010;
DRAM[37891] = 8'b10011011;
DRAM[37892] = 8'b10011100;
DRAM[37893] = 8'b10011100;
DRAM[37894] = 8'b10011101;
DRAM[37895] = 8'b10011101;
DRAM[37896] = 8'b10011100;
DRAM[37897] = 8'b10011100;
DRAM[37898] = 8'b10011101;
DRAM[37899] = 8'b10011110;
DRAM[37900] = 8'b10011110;
DRAM[37901] = 8'b10011111;
DRAM[37902] = 8'b10100000;
DRAM[37903] = 8'b10100000;
DRAM[37904] = 8'b10100001;
DRAM[37905] = 8'b10100001;
DRAM[37906] = 8'b10100000;
DRAM[37907] = 8'b10100000;
DRAM[37908] = 8'b10100001;
DRAM[37909] = 8'b10100001;
DRAM[37910] = 8'b10100010;
DRAM[37911] = 8'b10100011;
DRAM[37912] = 8'b10100101;
DRAM[37913] = 8'b10100100;
DRAM[37914] = 8'b10100011;
DRAM[37915] = 8'b10100011;
DRAM[37916] = 8'b10100010;
DRAM[37917] = 8'b10100011;
DRAM[37918] = 8'b10100011;
DRAM[37919] = 8'b10100100;
DRAM[37920] = 8'b10100100;
DRAM[37921] = 8'b10100101;
DRAM[37922] = 8'b10100101;
DRAM[37923] = 8'b10100110;
DRAM[37924] = 8'b10100110;
DRAM[37925] = 8'b10100101;
DRAM[37926] = 8'b10100100;
DRAM[37927] = 8'b10100100;
DRAM[37928] = 8'b10100101;
DRAM[37929] = 8'b10100100;
DRAM[37930] = 8'b10100100;
DRAM[37931] = 8'b10100011;
DRAM[37932] = 8'b10100011;
DRAM[37933] = 8'b10100100;
DRAM[37934] = 8'b10100100;
DRAM[37935] = 8'b10100101;
DRAM[37936] = 8'b10100110;
DRAM[37937] = 8'b10101011;
DRAM[37938] = 8'b10110001;
DRAM[37939] = 8'b10111000;
DRAM[37940] = 8'b11000010;
DRAM[37941] = 8'b11010010;
DRAM[37942] = 8'b11100100;
DRAM[37943] = 8'b11110001;
DRAM[37944] = 8'b11111010;
DRAM[37945] = 8'b11111001;
DRAM[37946] = 8'b11110111;
DRAM[37947] = 8'b11110111;
DRAM[37948] = 8'b11111010;
DRAM[37949] = 8'b11111011;
DRAM[37950] = 8'b11110011;
DRAM[37951] = 8'b11101001;
DRAM[37952] = 8'b11011010;
DRAM[37953] = 8'b11010100;
DRAM[37954] = 8'b11001100;
DRAM[37955] = 8'b11000101;
DRAM[37956] = 8'b11000001;
DRAM[37957] = 8'b10111100;
DRAM[37958] = 8'b10110101;
DRAM[37959] = 8'b10110000;
DRAM[37960] = 8'b10101110;
DRAM[37961] = 8'b10101110;
DRAM[37962] = 8'b10101101;
DRAM[37963] = 8'b10101010;
DRAM[37964] = 8'b10100111;
DRAM[37965] = 8'b10100110;
DRAM[37966] = 8'b10100111;
DRAM[37967] = 8'b10101000;
DRAM[37968] = 8'b10101100;
DRAM[37969] = 8'b10100110;
DRAM[37970] = 8'b10101111;
DRAM[37971] = 8'b10101110;
DRAM[37972] = 8'b10011100;
DRAM[37973] = 8'b10011111;
DRAM[37974] = 8'b10101100;
DRAM[37975] = 8'b10100111;
DRAM[37976] = 8'b10100111;
DRAM[37977] = 8'b10101011;
DRAM[37978] = 8'b10110000;
DRAM[37979] = 8'b10110011;
DRAM[37980] = 8'b10110011;
DRAM[37981] = 8'b10110011;
DRAM[37982] = 8'b10110101;
DRAM[37983] = 8'b10110111;
DRAM[37984] = 8'b10111111;
DRAM[37985] = 8'b11000100;
DRAM[37986] = 8'b11000101;
DRAM[37987] = 8'b10111110;
DRAM[37988] = 8'b10110101;
DRAM[37989] = 8'b10110111;
DRAM[37990] = 8'b11000111;
DRAM[37991] = 8'b11010110;
DRAM[37992] = 8'b11000111;
DRAM[37993] = 8'b11000010;
DRAM[37994] = 8'b11001001;
DRAM[37995] = 8'b11010001;
DRAM[37996] = 8'b11000001;
DRAM[37997] = 8'b10100111;
DRAM[37998] = 8'b10101000;
DRAM[37999] = 8'b10111110;
DRAM[38000] = 8'b10111010;
DRAM[38001] = 8'b11000011;
DRAM[38002] = 8'b11001010;
DRAM[38003] = 8'b11001000;
DRAM[38004] = 8'b11000111;
DRAM[38005] = 8'b11001111;
DRAM[38006] = 8'b11011011;
DRAM[38007] = 8'b11100100;
DRAM[38008] = 8'b11100000;
DRAM[38009] = 8'b11100101;
DRAM[38010] = 8'b11100110;
DRAM[38011] = 8'b11011111;
DRAM[38012] = 8'b11010100;
DRAM[38013] = 8'b11001110;
DRAM[38014] = 8'b11010010;
DRAM[38015] = 8'b11011000;
DRAM[38016] = 8'b11011010;
DRAM[38017] = 8'b11010000;
DRAM[38018] = 8'b11000100;
DRAM[38019] = 8'b10110011;
DRAM[38020] = 8'b10100111;
DRAM[38021] = 8'b10101000;
DRAM[38022] = 8'b10011110;
DRAM[38023] = 8'b10000101;
DRAM[38024] = 8'b1111111;
DRAM[38025] = 8'b1110100;
DRAM[38026] = 8'b1100110;
DRAM[38027] = 8'b1011101;
DRAM[38028] = 8'b1011100;
DRAM[38029] = 8'b1100001;
DRAM[38030] = 8'b1100111;
DRAM[38031] = 8'b1101100;
DRAM[38032] = 8'b1101101;
DRAM[38033] = 8'b1101100;
DRAM[38034] = 8'b1101010;
DRAM[38035] = 8'b1101001;
DRAM[38036] = 8'b1101010;
DRAM[38037] = 8'b1101100;
DRAM[38038] = 8'b1101110;
DRAM[38039] = 8'b1110000;
DRAM[38040] = 8'b1110111;
DRAM[38041] = 8'b10000001;
DRAM[38042] = 8'b1111110;
DRAM[38043] = 8'b1111010;
DRAM[38044] = 8'b1110111;
DRAM[38045] = 8'b1101001;
DRAM[38046] = 8'b1110110;
DRAM[38047] = 8'b10011111;
DRAM[38048] = 8'b10101101;
DRAM[38049] = 8'b11000001;
DRAM[38050] = 8'b11001111;
DRAM[38051] = 8'b11001111;
DRAM[38052] = 8'b11001111;
DRAM[38053] = 8'b11011011;
DRAM[38054] = 8'b11101000;
DRAM[38055] = 8'b11101110;
DRAM[38056] = 8'b11101100;
DRAM[38057] = 8'b11110010;
DRAM[38058] = 8'b11110011;
DRAM[38059] = 8'b11101110;
DRAM[38060] = 8'b11101110;
DRAM[38061] = 8'b11110010;
DRAM[38062] = 8'b11101110;
DRAM[38063] = 8'b11100110;
DRAM[38064] = 8'b11000110;
DRAM[38065] = 8'b10111010;
DRAM[38066] = 8'b10110010;
DRAM[38067] = 8'b10110111;
DRAM[38068] = 8'b10111111;
DRAM[38069] = 8'b11000001;
DRAM[38070] = 8'b10111111;
DRAM[38071] = 8'b10111110;
DRAM[38072] = 8'b10110111;
DRAM[38073] = 8'b10110010;
DRAM[38074] = 8'b10101111;
DRAM[38075] = 8'b10110001;
DRAM[38076] = 8'b10110110;
DRAM[38077] = 8'b10110111;
DRAM[38078] = 8'b10110100;
DRAM[38079] = 8'b10110001;
DRAM[38080] = 8'b10100111;
DRAM[38081] = 8'b10100101;
DRAM[38082] = 8'b10100111;
DRAM[38083] = 8'b10101110;
DRAM[38084] = 8'b10111000;
DRAM[38085] = 8'b11000111;
DRAM[38086] = 8'b11011011;
DRAM[38087] = 8'b11101101;
DRAM[38088] = 8'b11100111;
DRAM[38089] = 8'b11101001;
DRAM[38090] = 8'b11101110;
DRAM[38091] = 8'b11101000;
DRAM[38092] = 8'b11011000;
DRAM[38093] = 8'b11001110;
DRAM[38094] = 8'b10111111;
DRAM[38095] = 8'b10100110;
DRAM[38096] = 8'b10100001;
DRAM[38097] = 8'b10011011;
DRAM[38098] = 8'b10010110;
DRAM[38099] = 8'b10010101;
DRAM[38100] = 8'b10010100;
DRAM[38101] = 8'b10010000;
DRAM[38102] = 8'b10001110;
DRAM[38103] = 8'b10010000;
DRAM[38104] = 8'b10001111;
DRAM[38105] = 8'b10001110;
DRAM[38106] = 8'b10001101;
DRAM[38107] = 8'b10001101;
DRAM[38108] = 8'b10001100;
DRAM[38109] = 8'b10001100;
DRAM[38110] = 8'b10001101;
DRAM[38111] = 8'b10001101;
DRAM[38112] = 8'b10001011;
DRAM[38113] = 8'b10001011;
DRAM[38114] = 8'b10001010;
DRAM[38115] = 8'b10001001;
DRAM[38116] = 8'b10000111;
DRAM[38117] = 8'b10000101;
DRAM[38118] = 8'b10000011;
DRAM[38119] = 8'b10000001;
DRAM[38120] = 8'b10000001;
DRAM[38121] = 8'b10000001;
DRAM[38122] = 8'b10000000;
DRAM[38123] = 8'b1111111;
DRAM[38124] = 8'b1111111;
DRAM[38125] = 8'b1111111;
DRAM[38126] = 8'b1111111;
DRAM[38127] = 8'b10000000;
DRAM[38128] = 8'b1111111;
DRAM[38129] = 8'b1111110;
DRAM[38130] = 8'b1111101;
DRAM[38131] = 8'b1111100;
DRAM[38132] = 8'b1111011;
DRAM[38133] = 8'b1111100;
DRAM[38134] = 8'b1111101;
DRAM[38135] = 8'b1111110;
DRAM[38136] = 8'b1111100;
DRAM[38137] = 8'b1111100;
DRAM[38138] = 8'b1111100;
DRAM[38139] = 8'b1111100;
DRAM[38140] = 8'b1111100;
DRAM[38141] = 8'b1111100;
DRAM[38142] = 8'b1111100;
DRAM[38143] = 8'b1111100;
DRAM[38144] = 8'b10011010;
DRAM[38145] = 8'b10011010;
DRAM[38146] = 8'b10011010;
DRAM[38147] = 8'b10011011;
DRAM[38148] = 8'b10011100;
DRAM[38149] = 8'b10011101;
DRAM[38150] = 8'b10011101;
DRAM[38151] = 8'b10011110;
DRAM[38152] = 8'b10011011;
DRAM[38153] = 8'b10011100;
DRAM[38154] = 8'b10011100;
DRAM[38155] = 8'b10011101;
DRAM[38156] = 8'b10011111;
DRAM[38157] = 8'b10100000;
DRAM[38158] = 8'b10100000;
DRAM[38159] = 8'b10100001;
DRAM[38160] = 8'b10100001;
DRAM[38161] = 8'b10100001;
DRAM[38162] = 8'b10100001;
DRAM[38163] = 8'b10100001;
DRAM[38164] = 8'b10100001;
DRAM[38165] = 8'b10100010;
DRAM[38166] = 8'b10100011;
DRAM[38167] = 8'b10100011;
DRAM[38168] = 8'b10100101;
DRAM[38169] = 8'b10100100;
DRAM[38170] = 8'b10100100;
DRAM[38171] = 8'b10100011;
DRAM[38172] = 8'b10100011;
DRAM[38173] = 8'b10100100;
DRAM[38174] = 8'b10100101;
DRAM[38175] = 8'b10100101;
DRAM[38176] = 8'b10100110;
DRAM[38177] = 8'b10100110;
DRAM[38178] = 8'b10100110;
DRAM[38179] = 8'b10100111;
DRAM[38180] = 8'b10100110;
DRAM[38181] = 8'b10100101;
DRAM[38182] = 8'b10100100;
DRAM[38183] = 8'b10100100;
DRAM[38184] = 8'b10100101;
DRAM[38185] = 8'b10100100;
DRAM[38186] = 8'b10100100;
DRAM[38187] = 8'b10100011;
DRAM[38188] = 8'b10100011;
DRAM[38189] = 8'b10100100;
DRAM[38190] = 8'b10100100;
DRAM[38191] = 8'b10100101;
DRAM[38192] = 8'b10100111;
DRAM[38193] = 8'b10101011;
DRAM[38194] = 8'b10110100;
DRAM[38195] = 8'b11000001;
DRAM[38196] = 8'b11010001;
DRAM[38197] = 8'b11100010;
DRAM[38198] = 8'b11101111;
DRAM[38199] = 8'b11110111;
DRAM[38200] = 8'b11111010;
DRAM[38201] = 8'b11111011;
DRAM[38202] = 8'b11111011;
DRAM[38203] = 8'b11111010;
DRAM[38204] = 8'b11111100;
DRAM[38205] = 8'b11111100;
DRAM[38206] = 8'b11110100;
DRAM[38207] = 8'b11101001;
DRAM[38208] = 8'b11011010;
DRAM[38209] = 8'b11010100;
DRAM[38210] = 8'b11001011;
DRAM[38211] = 8'b11000101;
DRAM[38212] = 8'b11000000;
DRAM[38213] = 8'b10111011;
DRAM[38214] = 8'b10110100;
DRAM[38215] = 8'b10101111;
DRAM[38216] = 8'b10110001;
DRAM[38217] = 8'b10101111;
DRAM[38218] = 8'b10101101;
DRAM[38219] = 8'b10101010;
DRAM[38220] = 8'b10101000;
DRAM[38221] = 8'b10100110;
DRAM[38222] = 8'b10100101;
DRAM[38223] = 8'b10100100;
DRAM[38224] = 8'b10101101;
DRAM[38225] = 8'b10100101;
DRAM[38226] = 8'b10100010;
DRAM[38227] = 8'b10011101;
DRAM[38228] = 8'b10011000;
DRAM[38229] = 8'b10011101;
DRAM[38230] = 8'b10011111;
DRAM[38231] = 8'b10010110;
DRAM[38232] = 8'b10011110;
DRAM[38233] = 8'b10100000;
DRAM[38234] = 8'b10100011;
DRAM[38235] = 8'b10101011;
DRAM[38236] = 8'b10110100;
DRAM[38237] = 8'b10111100;
DRAM[38238] = 8'b11000000;
DRAM[38239] = 8'b11000001;
DRAM[38240] = 8'b10111011;
DRAM[38241] = 8'b11000010;
DRAM[38242] = 8'b11001000;
DRAM[38243] = 8'b11000111;
DRAM[38244] = 8'b11000011;
DRAM[38245] = 8'b11000100;
DRAM[38246] = 8'b11001100;
DRAM[38247] = 8'b11010101;
DRAM[38248] = 8'b11001001;
DRAM[38249] = 8'b11000111;
DRAM[38250] = 8'b11000001;
DRAM[38251] = 8'b10111000;
DRAM[38252] = 8'b10110000;
DRAM[38253] = 8'b10101101;
DRAM[38254] = 8'b10110011;
DRAM[38255] = 8'b10111010;
DRAM[38256] = 8'b11000010;
DRAM[38257] = 8'b11000100;
DRAM[38258] = 8'b11000110;
DRAM[38259] = 8'b11000101;
DRAM[38260] = 8'b11000110;
DRAM[38261] = 8'b11001110;
DRAM[38262] = 8'b11011011;
DRAM[38263] = 8'b11100101;
DRAM[38264] = 8'b11011000;
DRAM[38265] = 8'b11011101;
DRAM[38266] = 8'b11100011;
DRAM[38267] = 8'b11100110;
DRAM[38268] = 8'b11100101;
DRAM[38269] = 8'b11100100;
DRAM[38270] = 8'b11100101;
DRAM[38271] = 8'b11100111;
DRAM[38272] = 8'b11100000;
DRAM[38273] = 8'b11011101;
DRAM[38274] = 8'b11010011;
DRAM[38275] = 8'b10111110;
DRAM[38276] = 8'b10101101;
DRAM[38277] = 8'b10101010;
DRAM[38278] = 8'b10011001;
DRAM[38279] = 8'b1110111;
DRAM[38280] = 8'b1100100;
DRAM[38281] = 8'b1100010;
DRAM[38282] = 8'b1011111;
DRAM[38283] = 8'b1011011;
DRAM[38284] = 8'b1011010;
DRAM[38285] = 8'b1011110;
DRAM[38286] = 8'b1100101;
DRAM[38287] = 8'b1101011;
DRAM[38288] = 8'b1110111;
DRAM[38289] = 8'b1110110;
DRAM[38290] = 8'b1110100;
DRAM[38291] = 8'b1110001;
DRAM[38292] = 8'b1110000;
DRAM[38293] = 8'b1101111;
DRAM[38294] = 8'b1101111;
DRAM[38295] = 8'b1110000;
DRAM[38296] = 8'b1111100;
DRAM[38297] = 8'b10000010;
DRAM[38298] = 8'b10000100;
DRAM[38299] = 8'b10001000;
DRAM[38300] = 8'b10001100;
DRAM[38301] = 8'b10000010;
DRAM[38302] = 8'b1110110;
DRAM[38303] = 8'b1110111;
DRAM[38304] = 8'b10011101;
DRAM[38305] = 8'b10110101;
DRAM[38306] = 8'b11000100;
DRAM[38307] = 8'b10111111;
DRAM[38308] = 8'b10111100;
DRAM[38309] = 8'b11001001;
DRAM[38310] = 8'b11011000;
DRAM[38311] = 8'b11011111;
DRAM[38312] = 8'b11011111;
DRAM[38313] = 8'b11101011;
DRAM[38314] = 8'b11110000;
DRAM[38315] = 8'b11101101;
DRAM[38316] = 8'b11101100;
DRAM[38317] = 8'b11110010;
DRAM[38318] = 8'b11110100;
DRAM[38319] = 8'b11110000;
DRAM[38320] = 8'b11100111;
DRAM[38321] = 8'b11001111;
DRAM[38322] = 8'b10111011;
DRAM[38323] = 8'b10111001;
DRAM[38324] = 8'b10111111;
DRAM[38325] = 8'b10111111;
DRAM[38326] = 8'b10111110;
DRAM[38327] = 8'b10111111;
DRAM[38328] = 8'b10110111;
DRAM[38329] = 8'b10110001;
DRAM[38330] = 8'b10101110;
DRAM[38331] = 8'b10110011;
DRAM[38332] = 8'b10111000;
DRAM[38333] = 8'b10110110;
DRAM[38334] = 8'b10110010;
DRAM[38335] = 8'b10110000;
DRAM[38336] = 8'b10101001;
DRAM[38337] = 8'b10100111;
DRAM[38338] = 8'b10101010;
DRAM[38339] = 8'b10110011;
DRAM[38340] = 8'b10111111;
DRAM[38341] = 8'b11001100;
DRAM[38342] = 8'b11011101;
DRAM[38343] = 8'b11101100;
DRAM[38344] = 8'b11101101;
DRAM[38345] = 8'b11101111;
DRAM[38346] = 8'b11110110;
DRAM[38347] = 8'b11110010;
DRAM[38348] = 8'b11100110;
DRAM[38349] = 8'b11100010;
DRAM[38350] = 8'b11011000;
DRAM[38351] = 8'b11000010;
DRAM[38352] = 8'b10101001;
DRAM[38353] = 8'b10100010;
DRAM[38354] = 8'b10011100;
DRAM[38355] = 8'b10011010;
DRAM[38356] = 8'b10010111;
DRAM[38357] = 8'b10010001;
DRAM[38358] = 8'b10001101;
DRAM[38359] = 8'b10001110;
DRAM[38360] = 8'b10001111;
DRAM[38361] = 8'b10001111;
DRAM[38362] = 8'b10001110;
DRAM[38363] = 8'b10001101;
DRAM[38364] = 8'b10001101;
DRAM[38365] = 8'b10001101;
DRAM[38366] = 8'b10001101;
DRAM[38367] = 8'b10001101;
DRAM[38368] = 8'b10001010;
DRAM[38369] = 8'b10001010;
DRAM[38370] = 8'b10001001;
DRAM[38371] = 8'b10001001;
DRAM[38372] = 8'b10000111;
DRAM[38373] = 8'b10000101;
DRAM[38374] = 8'b10000011;
DRAM[38375] = 8'b10000010;
DRAM[38376] = 8'b10000001;
DRAM[38377] = 8'b10000000;
DRAM[38378] = 8'b10000000;
DRAM[38379] = 8'b1111111;
DRAM[38380] = 8'b1111111;
DRAM[38381] = 8'b1111111;
DRAM[38382] = 8'b10000000;
DRAM[38383] = 8'b10000001;
DRAM[38384] = 8'b1111111;
DRAM[38385] = 8'b1111110;
DRAM[38386] = 8'b1111100;
DRAM[38387] = 8'b1111011;
DRAM[38388] = 8'b1111011;
DRAM[38389] = 8'b1111100;
DRAM[38390] = 8'b1111101;
DRAM[38391] = 8'b1111110;
DRAM[38392] = 8'b1111101;
DRAM[38393] = 8'b1111101;
DRAM[38394] = 8'b1111101;
DRAM[38395] = 8'b1111101;
DRAM[38396] = 8'b1111101;
DRAM[38397] = 8'b1111101;
DRAM[38398] = 8'b1111101;
DRAM[38399] = 8'b1111101;
DRAM[38400] = 8'b10011010;
DRAM[38401] = 8'b10011010;
DRAM[38402] = 8'b10011011;
DRAM[38403] = 8'b10011011;
DRAM[38404] = 8'b10011100;
DRAM[38405] = 8'b10011101;
DRAM[38406] = 8'b10011110;
DRAM[38407] = 8'b10011110;
DRAM[38408] = 8'b10011011;
DRAM[38409] = 8'b10011011;
DRAM[38410] = 8'b10011100;
DRAM[38411] = 8'b10011101;
DRAM[38412] = 8'b10011111;
DRAM[38413] = 8'b10100000;
DRAM[38414] = 8'b10100001;
DRAM[38415] = 8'b10100001;
DRAM[38416] = 8'b10100010;
DRAM[38417] = 8'b10100001;
DRAM[38418] = 8'b10100001;
DRAM[38419] = 8'b10100001;
DRAM[38420] = 8'b10100001;
DRAM[38421] = 8'b10100010;
DRAM[38422] = 8'b10100011;
DRAM[38423] = 8'b10100100;
DRAM[38424] = 8'b10100100;
DRAM[38425] = 8'b10100100;
DRAM[38426] = 8'b10100011;
DRAM[38427] = 8'b10100100;
DRAM[38428] = 8'b10100100;
DRAM[38429] = 8'b10100101;
DRAM[38430] = 8'b10100111;
DRAM[38431] = 8'b10100111;
DRAM[38432] = 8'b10100111;
DRAM[38433] = 8'b10100111;
DRAM[38434] = 8'b10100111;
DRAM[38435] = 8'b10101000;
DRAM[38436] = 8'b10100111;
DRAM[38437] = 8'b10100110;
DRAM[38438] = 8'b10100101;
DRAM[38439] = 8'b10100100;
DRAM[38440] = 8'b10100101;
DRAM[38441] = 8'b10100100;
DRAM[38442] = 8'b10100100;
DRAM[38443] = 8'b10100011;
DRAM[38444] = 8'b10100011;
DRAM[38445] = 8'b10100100;
DRAM[38446] = 8'b10100100;
DRAM[38447] = 8'b10100101;
DRAM[38448] = 8'b10101100;
DRAM[38449] = 8'b10101101;
DRAM[38450] = 8'b10110100;
DRAM[38451] = 8'b11000110;
DRAM[38452] = 8'b11011101;
DRAM[38453] = 8'b11110010;
DRAM[38454] = 8'b11111111;
DRAM[38455] = 8'b11111111;
DRAM[38456] = 8'b11111100;
DRAM[38457] = 8'b11111110;
DRAM[38458] = 8'b11111111;
DRAM[38459] = 8'b11111101;
DRAM[38460] = 8'b11111110;
DRAM[38461] = 8'b11111101;
DRAM[38462] = 8'b11110110;
DRAM[38463] = 8'b11101110;
DRAM[38464] = 8'b11100010;
DRAM[38465] = 8'b11011001;
DRAM[38466] = 8'b11001110;
DRAM[38467] = 8'b11000101;
DRAM[38468] = 8'b11000000;
DRAM[38469] = 8'b10111100;
DRAM[38470] = 8'b10111000;
DRAM[38471] = 8'b10110100;
DRAM[38472] = 8'b10110110;
DRAM[38473] = 8'b10110011;
DRAM[38474] = 8'b10101111;
DRAM[38475] = 8'b10101110;
DRAM[38476] = 8'b10101110;
DRAM[38477] = 8'b10101100;
DRAM[38478] = 8'b10101000;
DRAM[38479] = 8'b10100101;
DRAM[38480] = 8'b10011100;
DRAM[38481] = 8'b10100001;
DRAM[38482] = 8'b10011100;
DRAM[38483] = 8'b10011011;
DRAM[38484] = 8'b10100111;
DRAM[38485] = 8'b10101111;
DRAM[38486] = 8'b10101101;
DRAM[38487] = 8'b10101011;
DRAM[38488] = 8'b10011011;
DRAM[38489] = 8'b10011000;
DRAM[38490] = 8'b10011010;
DRAM[38491] = 8'b10100100;
DRAM[38492] = 8'b10110100;
DRAM[38493] = 8'b11000001;
DRAM[38494] = 8'b11000110;
DRAM[38495] = 8'b11000101;
DRAM[38496] = 8'b10111101;
DRAM[38497] = 8'b10111101;
DRAM[38498] = 8'b11000000;
DRAM[38499] = 8'b11001000;
DRAM[38500] = 8'b11010000;
DRAM[38501] = 8'b11010000;
DRAM[38502] = 8'b11001001;
DRAM[38503] = 8'b11000001;
DRAM[38504] = 8'b11000011;
DRAM[38505] = 8'b10111111;
DRAM[38506] = 8'b10110011;
DRAM[38507] = 8'b10101001;
DRAM[38508] = 8'b10110000;
DRAM[38509] = 8'b10111111;
DRAM[38510] = 8'b10111111;
DRAM[38511] = 8'b10110101;
DRAM[38512] = 8'b11001000;
DRAM[38513] = 8'b11001000;
DRAM[38514] = 8'b11001001;
DRAM[38515] = 8'b11001011;
DRAM[38516] = 8'b11001111;
DRAM[38517] = 8'b11010100;
DRAM[38518] = 8'b11011011;
DRAM[38519] = 8'b11100001;
DRAM[38520] = 8'b11010111;
DRAM[38521] = 8'b11011010;
DRAM[38522] = 8'b11100001;
DRAM[38523] = 8'b11101011;
DRAM[38524] = 8'b11110011;
DRAM[38525] = 8'b11110011;
DRAM[38526] = 8'b11101110;
DRAM[38527] = 8'b11101000;
DRAM[38528] = 8'b11010111;
DRAM[38529] = 8'b11001111;
DRAM[38530] = 8'b11001011;
DRAM[38531] = 8'b11000110;
DRAM[38532] = 8'b10111010;
DRAM[38533] = 8'b10101100;
DRAM[38534] = 8'b10010000;
DRAM[38535] = 8'b1101101;
DRAM[38536] = 8'b1011000;
DRAM[38537] = 8'b1011111;
DRAM[38538] = 8'b1100100;
DRAM[38539] = 8'b1100011;
DRAM[38540] = 8'b1011110;
DRAM[38541] = 8'b1011101;
DRAM[38542] = 8'b1100010;
DRAM[38543] = 8'b1100111;
DRAM[38544] = 8'b1110101;
DRAM[38545] = 8'b1110100;
DRAM[38546] = 8'b1110011;
DRAM[38547] = 8'b1110010;
DRAM[38548] = 8'b1110001;
DRAM[38549] = 8'b1110000;
DRAM[38550] = 8'b1110000;
DRAM[38551] = 8'b1110000;
DRAM[38552] = 8'b1111010;
DRAM[38553] = 8'b1111010;
DRAM[38554] = 8'b1111111;
DRAM[38555] = 8'b10000111;
DRAM[38556] = 8'b10010010;
DRAM[38557] = 8'b10011110;
DRAM[38558] = 8'b10010001;
DRAM[38559] = 8'b1110011;
DRAM[38560] = 8'b10000100;
DRAM[38561] = 8'b10100001;
DRAM[38562] = 8'b10110110;
DRAM[38563] = 8'b10110010;
DRAM[38564] = 8'b10101110;
DRAM[38565] = 8'b10111010;
DRAM[38566] = 8'b11001010;
DRAM[38567] = 8'b11010000;
DRAM[38568] = 8'b11010111;
DRAM[38569] = 8'b11100110;
DRAM[38570] = 8'b11110000;
DRAM[38571] = 8'b11101101;
DRAM[38572] = 8'b11101010;
DRAM[38573] = 8'b11110000;
DRAM[38574] = 8'b11110101;
DRAM[38575] = 8'b11110100;
DRAM[38576] = 8'b11100011;
DRAM[38577] = 8'b11001101;
DRAM[38578] = 8'b10111100;
DRAM[38579] = 8'b10111100;
DRAM[38580] = 8'b11000010;
DRAM[38581] = 8'b11000100;
DRAM[38582] = 8'b11000111;
DRAM[38583] = 8'b11001101;
DRAM[38584] = 8'b11000000;
DRAM[38585] = 8'b10110111;
DRAM[38586] = 8'b10110010;
DRAM[38587] = 8'b10110110;
DRAM[38588] = 8'b10111001;
DRAM[38589] = 8'b10110110;
DRAM[38590] = 8'b10110010;
DRAM[38591] = 8'b10110001;
DRAM[38592] = 8'b10101110;
DRAM[38593] = 8'b10101011;
DRAM[38594] = 8'b10101101;
DRAM[38595] = 8'b10111000;
DRAM[38596] = 8'b11000100;
DRAM[38597] = 8'b11001111;
DRAM[38598] = 8'b11011010;
DRAM[38599] = 8'b11100011;
DRAM[38600] = 8'b11110000;
DRAM[38601] = 8'b11101110;
DRAM[38602] = 8'b11101110;
DRAM[38603] = 8'b11100110;
DRAM[38604] = 8'b11011011;
DRAM[38605] = 8'b11011101;
DRAM[38606] = 8'b11011001;
DRAM[38607] = 8'b11001001;
DRAM[38608] = 8'b10100111;
DRAM[38609] = 8'b10100000;
DRAM[38610] = 8'b10011011;
DRAM[38611] = 8'b10011010;
DRAM[38612] = 8'b10010111;
DRAM[38613] = 8'b10010010;
DRAM[38614] = 8'b10001110;
DRAM[38615] = 8'b10001111;
DRAM[38616] = 8'b10010000;
DRAM[38617] = 8'b10001111;
DRAM[38618] = 8'b10001110;
DRAM[38619] = 8'b10001101;
DRAM[38620] = 8'b10001101;
DRAM[38621] = 8'b10001101;
DRAM[38622] = 8'b10001101;
DRAM[38623] = 8'b10001110;
DRAM[38624] = 8'b10001001;
DRAM[38625] = 8'b10001001;
DRAM[38626] = 8'b10001001;
DRAM[38627] = 8'b10001000;
DRAM[38628] = 8'b10000111;
DRAM[38629] = 8'b10000110;
DRAM[38630] = 8'b10000101;
DRAM[38631] = 8'b10000100;
DRAM[38632] = 8'b10000001;
DRAM[38633] = 8'b10000001;
DRAM[38634] = 8'b10000000;
DRAM[38635] = 8'b10000000;
DRAM[38636] = 8'b10000000;
DRAM[38637] = 8'b10000000;
DRAM[38638] = 8'b10000001;
DRAM[38639] = 8'b10000010;
DRAM[38640] = 8'b1111110;
DRAM[38641] = 8'b1111110;
DRAM[38642] = 8'b1111100;
DRAM[38643] = 8'b1111011;
DRAM[38644] = 8'b1111011;
DRAM[38645] = 8'b1111100;
DRAM[38646] = 8'b1111110;
DRAM[38647] = 8'b1111111;
DRAM[38648] = 8'b1111101;
DRAM[38649] = 8'b1111101;
DRAM[38650] = 8'b1111101;
DRAM[38651] = 8'b1111101;
DRAM[38652] = 8'b1111101;
DRAM[38653] = 8'b1111101;
DRAM[38654] = 8'b1111101;
DRAM[38655] = 8'b1111101;
DRAM[38656] = 8'b10011010;
DRAM[38657] = 8'b10011010;
DRAM[38658] = 8'b10011011;
DRAM[38659] = 8'b10011100;
DRAM[38660] = 8'b10011100;
DRAM[38661] = 8'b10011101;
DRAM[38662] = 8'b10011110;
DRAM[38663] = 8'b10011110;
DRAM[38664] = 8'b10011010;
DRAM[38665] = 8'b10011011;
DRAM[38666] = 8'b10011100;
DRAM[38667] = 8'b10011101;
DRAM[38668] = 8'b10011111;
DRAM[38669] = 8'b10100000;
DRAM[38670] = 8'b10100001;
DRAM[38671] = 8'b10100010;
DRAM[38672] = 8'b10100010;
DRAM[38673] = 8'b10100001;
DRAM[38674] = 8'b10100001;
DRAM[38675] = 8'b10100001;
DRAM[38676] = 8'b10100001;
DRAM[38677] = 8'b10100010;
DRAM[38678] = 8'b10100011;
DRAM[38679] = 8'b10100100;
DRAM[38680] = 8'b10100011;
DRAM[38681] = 8'b10100011;
DRAM[38682] = 8'b10100011;
DRAM[38683] = 8'b10100100;
DRAM[38684] = 8'b10100101;
DRAM[38685] = 8'b10100110;
DRAM[38686] = 8'b10101000;
DRAM[38687] = 8'b10101001;
DRAM[38688] = 8'b10101000;
DRAM[38689] = 8'b10101000;
DRAM[38690] = 8'b10101000;
DRAM[38691] = 8'b10101000;
DRAM[38692] = 8'b10101000;
DRAM[38693] = 8'b10100111;
DRAM[38694] = 8'b10100110;
DRAM[38695] = 8'b10100101;
DRAM[38696] = 8'b10100101;
DRAM[38697] = 8'b10100100;
DRAM[38698] = 8'b10100100;
DRAM[38699] = 8'b10100011;
DRAM[38700] = 8'b10100011;
DRAM[38701] = 8'b10100100;
DRAM[38702] = 8'b10100100;
DRAM[38703] = 8'b10100101;
DRAM[38704] = 8'b10101011;
DRAM[38705] = 8'b10110001;
DRAM[38706] = 8'b11000000;
DRAM[38707] = 8'b11011001;
DRAM[38708] = 8'b11110001;
DRAM[38709] = 8'b11111110;
DRAM[38710] = 8'b11111101;
DRAM[38711] = 8'b11110111;
DRAM[38712] = 8'b11111011;
DRAM[38713] = 8'b11111110;
DRAM[38714] = 8'b11111111;
DRAM[38715] = 8'b11111101;
DRAM[38716] = 8'b11111110;
DRAM[38717] = 8'b11111110;
DRAM[38718] = 8'b11111010;
DRAM[38719] = 8'b11110100;
DRAM[38720] = 8'b11101011;
DRAM[38721] = 8'b11100000;
DRAM[38722] = 8'b11010001;
DRAM[38723] = 8'b11000110;
DRAM[38724] = 8'b11000001;
DRAM[38725] = 8'b10111111;
DRAM[38726] = 8'b10111110;
DRAM[38727] = 8'b10111100;
DRAM[38728] = 8'b10110111;
DRAM[38729] = 8'b10110010;
DRAM[38730] = 8'b10101110;
DRAM[38731] = 8'b10101110;
DRAM[38732] = 8'b10110000;
DRAM[38733] = 8'b10101111;
DRAM[38734] = 8'b10101001;
DRAM[38735] = 8'b10100011;
DRAM[38736] = 8'b10100000;
DRAM[38737] = 8'b10110001;
DRAM[38738] = 8'b10101001;
DRAM[38739] = 8'b10011010;
DRAM[38740] = 8'b10011011;
DRAM[38741] = 8'b10010100;
DRAM[38742] = 8'b10001010;
DRAM[38743] = 8'b10010000;
DRAM[38744] = 8'b10100000;
DRAM[38745] = 8'b10100001;
DRAM[38746] = 8'b10101001;
DRAM[38747] = 8'b10111001;
DRAM[38748] = 8'b11000110;
DRAM[38749] = 8'b11000110;
DRAM[38750] = 8'b10111001;
DRAM[38751] = 8'b10101011;
DRAM[38752] = 8'b10111001;
DRAM[38753] = 8'b11000001;
DRAM[38754] = 8'b11001100;
DRAM[38755] = 8'b11010000;
DRAM[38756] = 8'b11001101;
DRAM[38757] = 8'b11000111;
DRAM[38758] = 8'b11000101;
DRAM[38759] = 8'b11000101;
DRAM[38760] = 8'b10110010;
DRAM[38761] = 8'b10111000;
DRAM[38762] = 8'b10111101;
DRAM[38763] = 8'b10111110;
DRAM[38764] = 8'b10111101;
DRAM[38765] = 8'b11000000;
DRAM[38766] = 8'b11000110;
DRAM[38767] = 8'b11001011;
DRAM[38768] = 8'b10111100;
DRAM[38769] = 8'b10111101;
DRAM[38770] = 8'b11000011;
DRAM[38771] = 8'b11001101;
DRAM[38772] = 8'b11010111;
DRAM[38773] = 8'b11011100;
DRAM[38774] = 8'b11100001;
DRAM[38775] = 8'b11100100;
DRAM[38776] = 8'b11101001;
DRAM[38777] = 8'b11100111;
DRAM[38778] = 8'b11101001;
DRAM[38779] = 8'b11110000;
DRAM[38780] = 8'b11110101;
DRAM[38781] = 8'b11101111;
DRAM[38782] = 8'b11100000;
DRAM[38783] = 8'b11010010;
DRAM[38784] = 8'b11001101;
DRAM[38785] = 8'b10111011;
DRAM[38786] = 8'b10111001;
DRAM[38787] = 8'b11000001;
DRAM[38788] = 8'b10111000;
DRAM[38789] = 8'b10011101;
DRAM[38790] = 8'b1110110;
DRAM[38791] = 8'b1010011;
DRAM[38792] = 8'b1011010;
DRAM[38793] = 8'b1100101;
DRAM[38794] = 8'b1101111;
DRAM[38795] = 8'b1101111;
DRAM[38796] = 8'b1100110;
DRAM[38797] = 8'b1100000;
DRAM[38798] = 8'b1100001;
DRAM[38799] = 8'b1100110;
DRAM[38800] = 8'b1100101;
DRAM[38801] = 8'b1100110;
DRAM[38802] = 8'b1100110;
DRAM[38803] = 8'b1101000;
DRAM[38804] = 8'b1101001;
DRAM[38805] = 8'b1101010;
DRAM[38806] = 8'b1101011;
DRAM[38807] = 8'b1101100;
DRAM[38808] = 8'b1110001;
DRAM[38809] = 8'b1101110;
DRAM[38810] = 8'b1110011;
DRAM[38811] = 8'b1110101;
DRAM[38812] = 8'b10000001;
DRAM[38813] = 8'b10100100;
DRAM[38814] = 8'b10101011;
DRAM[38815] = 8'b10001001;
DRAM[38816] = 8'b1011110;
DRAM[38817] = 8'b10000010;
DRAM[38818] = 8'b10011111;
DRAM[38819] = 8'b10100010;
DRAM[38820] = 8'b10100100;
DRAM[38821] = 8'b10110101;
DRAM[38822] = 8'b11001000;
DRAM[38823] = 8'b11001111;
DRAM[38824] = 8'b11010101;
DRAM[38825] = 8'b11100110;
DRAM[38826] = 8'b11110000;
DRAM[38827] = 8'b11101100;
DRAM[38828] = 8'b11101000;
DRAM[38829] = 8'b11101011;
DRAM[38830] = 8'b11110000;
DRAM[38831] = 8'b11110001;
DRAM[38832] = 8'b11100101;
DRAM[38833] = 8'b11010011;
DRAM[38834] = 8'b11000101;
DRAM[38835] = 8'b11000010;
DRAM[38836] = 8'b10111101;
DRAM[38837] = 8'b10110011;
DRAM[38838] = 8'b10101111;
DRAM[38839] = 8'b10110011;
DRAM[38840] = 8'b11001001;
DRAM[38841] = 8'b10111110;
DRAM[38842] = 8'b10110110;
DRAM[38843] = 8'b10111000;
DRAM[38844] = 8'b10111001;
DRAM[38845] = 8'b10110110;
DRAM[38846] = 8'b10110010;
DRAM[38847] = 8'b10110011;
DRAM[38848] = 8'b10101111;
DRAM[38849] = 8'b10101100;
DRAM[38850] = 8'b10110000;
DRAM[38851] = 8'b10111110;
DRAM[38852] = 8'b11001110;
DRAM[38853] = 8'b11011001;
DRAM[38854] = 8'b11100011;
DRAM[38855] = 8'b11101010;
DRAM[38856] = 8'b11101010;
DRAM[38857] = 8'b11101011;
DRAM[38858] = 8'b11101101;
DRAM[38859] = 8'b11100100;
DRAM[38860] = 8'b11010011;
DRAM[38861] = 8'b11001001;
DRAM[38862] = 8'b10111010;
DRAM[38863] = 8'b10100010;
DRAM[38864] = 8'b10011101;
DRAM[38865] = 8'b10010111;
DRAM[38866] = 8'b10010100;
DRAM[38867] = 8'b10010110;
DRAM[38868] = 8'b10010101;
DRAM[38869] = 8'b10010010;
DRAM[38870] = 8'b10010000;
DRAM[38871] = 8'b10010010;
DRAM[38872] = 8'b10010000;
DRAM[38873] = 8'b10001111;
DRAM[38874] = 8'b10001110;
DRAM[38875] = 8'b10001101;
DRAM[38876] = 8'b10001101;
DRAM[38877] = 8'b10001101;
DRAM[38878] = 8'b10001101;
DRAM[38879] = 8'b10001110;
DRAM[38880] = 8'b10001000;
DRAM[38881] = 8'b10001000;
DRAM[38882] = 8'b10001000;
DRAM[38883] = 8'b10001000;
DRAM[38884] = 8'b10001000;
DRAM[38885] = 8'b10000110;
DRAM[38886] = 8'b10000101;
DRAM[38887] = 8'b10000101;
DRAM[38888] = 8'b10000010;
DRAM[38889] = 8'b10000001;
DRAM[38890] = 8'b10000001;
DRAM[38891] = 8'b10000000;
DRAM[38892] = 8'b10000000;
DRAM[38893] = 8'b10000001;
DRAM[38894] = 8'b10000010;
DRAM[38895] = 8'b10000010;
DRAM[38896] = 8'b1111110;
DRAM[38897] = 8'b1111101;
DRAM[38898] = 8'b1111100;
DRAM[38899] = 8'b1111011;
DRAM[38900] = 8'b1111011;
DRAM[38901] = 8'b1111101;
DRAM[38902] = 8'b1111110;
DRAM[38903] = 8'b1111111;
DRAM[38904] = 8'b1111101;
DRAM[38905] = 8'b1111101;
DRAM[38906] = 8'b1111101;
DRAM[38907] = 8'b1111101;
DRAM[38908] = 8'b1111101;
DRAM[38909] = 8'b1111101;
DRAM[38910] = 8'b1111101;
DRAM[38911] = 8'b1111101;
DRAM[38912] = 8'b10011010;
DRAM[38913] = 8'b10011010;
DRAM[38914] = 8'b10011010;
DRAM[38915] = 8'b10011011;
DRAM[38916] = 8'b10011011;
DRAM[38917] = 8'b10011100;
DRAM[38918] = 8'b10011100;
DRAM[38919] = 8'b10011100;
DRAM[38920] = 8'b10011100;
DRAM[38921] = 8'b10011100;
DRAM[38922] = 8'b10011100;
DRAM[38923] = 8'b10011101;
DRAM[38924] = 8'b10011110;
DRAM[38925] = 8'b10011111;
DRAM[38926] = 8'b10100001;
DRAM[38927] = 8'b10100001;
DRAM[38928] = 8'b10100001;
DRAM[38929] = 8'b10100001;
DRAM[38930] = 8'b10100010;
DRAM[38931] = 8'b10100011;
DRAM[38932] = 8'b10100011;
DRAM[38933] = 8'b10100100;
DRAM[38934] = 8'b10100101;
DRAM[38935] = 8'b10100101;
DRAM[38936] = 8'b10100101;
DRAM[38937] = 8'b10100100;
DRAM[38938] = 8'b10100100;
DRAM[38939] = 8'b10100100;
DRAM[38940] = 8'b10100100;
DRAM[38941] = 8'b10100101;
DRAM[38942] = 8'b10100110;
DRAM[38943] = 8'b10100111;
DRAM[38944] = 8'b10101000;
DRAM[38945] = 8'b10101000;
DRAM[38946] = 8'b10100111;
DRAM[38947] = 8'b10100110;
DRAM[38948] = 8'b10100110;
DRAM[38949] = 8'b10100101;
DRAM[38950] = 8'b10100100;
DRAM[38951] = 8'b10100100;
DRAM[38952] = 8'b10100110;
DRAM[38953] = 8'b10100011;
DRAM[38954] = 8'b10100010;
DRAM[38955] = 8'b10100100;
DRAM[38956] = 8'b10100100;
DRAM[38957] = 8'b10100010;
DRAM[38958] = 8'b10100100;
DRAM[38959] = 8'b10101001;
DRAM[38960] = 8'b10110001;
DRAM[38961] = 8'b10111100;
DRAM[38962] = 8'b11010011;
DRAM[38963] = 8'b11101101;
DRAM[38964] = 8'b11111011;
DRAM[38965] = 8'b11111101;
DRAM[38966] = 8'b11111101;
DRAM[38967] = 8'b11111111;
DRAM[38968] = 8'b11111101;
DRAM[38969] = 8'b11111100;
DRAM[38970] = 8'b11111100;
DRAM[38971] = 8'b11111101;
DRAM[38972] = 8'b11111110;
DRAM[38973] = 8'b11111100;
DRAM[38974] = 8'b11111000;
DRAM[38975] = 8'b11110100;
DRAM[38976] = 8'b11101010;
DRAM[38977] = 8'b11011110;
DRAM[38978] = 8'b11001111;
DRAM[38979] = 8'b11000101;
DRAM[38980] = 8'b11000000;
DRAM[38981] = 8'b10111011;
DRAM[38982] = 8'b10110011;
DRAM[38983] = 8'b10101011;
DRAM[38984] = 8'b10100011;
DRAM[38985] = 8'b10100111;
DRAM[38986] = 8'b10101000;
DRAM[38987] = 8'b10100110;
DRAM[38988] = 8'b10101000;
DRAM[38989] = 8'b10101100;
DRAM[38990] = 8'b10101010;
DRAM[38991] = 8'b10100011;
DRAM[38992] = 8'b10100101;
DRAM[38993] = 8'b10011011;
DRAM[38994] = 8'b10010011;
DRAM[38995] = 8'b10010011;
DRAM[38996] = 8'b10010111;
DRAM[38997] = 8'b10011011;
DRAM[38998] = 8'b10100010;
DRAM[38999] = 8'b10101001;
DRAM[39000] = 8'b10101101;
DRAM[39001] = 8'b10111001;
DRAM[39002] = 8'b11000000;
DRAM[39003] = 8'b10111001;
DRAM[39004] = 8'b10110100;
DRAM[39005] = 8'b10111000;
DRAM[39006] = 8'b11000001;
DRAM[39007] = 8'b11000110;
DRAM[39008] = 8'b11000111;
DRAM[39009] = 8'b11000100;
DRAM[39010] = 8'b10111110;
DRAM[39011] = 8'b10110111;
DRAM[39012] = 8'b10110010;
DRAM[39013] = 8'b10110010;
DRAM[39014] = 8'b10110111;
DRAM[39015] = 8'b10111100;
DRAM[39016] = 8'b10111000;
DRAM[39017] = 8'b10111111;
DRAM[39018] = 8'b11000110;
DRAM[39019] = 8'b11000100;
DRAM[39020] = 8'b10111100;
DRAM[39021] = 8'b10111001;
DRAM[39022] = 8'b10111111;
DRAM[39023] = 8'b11000111;
DRAM[39024] = 8'b10110001;
DRAM[39025] = 8'b10110111;
DRAM[39026] = 8'b11000111;
DRAM[39027] = 8'b11010111;
DRAM[39028] = 8'b11011010;
DRAM[39029] = 8'b11010101;
DRAM[39030] = 8'b11011010;
DRAM[39031] = 8'b11100101;
DRAM[39032] = 8'b11100001;
DRAM[39033] = 8'b11011101;
DRAM[39034] = 8'b11101010;
DRAM[39035] = 8'b11110001;
DRAM[39036] = 8'b11100111;
DRAM[39037] = 8'b11100111;
DRAM[39038] = 8'b11100010;
DRAM[39039] = 8'b11001011;
DRAM[39040] = 8'b11000100;
DRAM[39041] = 8'b11010100;
DRAM[39042] = 8'b10111100;
DRAM[39043] = 8'b10101111;
DRAM[39044] = 8'b10100100;
DRAM[39045] = 8'b1111101;
DRAM[39046] = 8'b1100011;
DRAM[39047] = 8'b1010111;
DRAM[39048] = 8'b1110011;
DRAM[39049] = 8'b1111011;
DRAM[39050] = 8'b1111110;
DRAM[39051] = 8'b1110111;
DRAM[39052] = 8'b1101010;
DRAM[39053] = 8'b1100001;
DRAM[39054] = 8'b1011111;
DRAM[39055] = 8'b1100000;
DRAM[39056] = 8'b1011010;
DRAM[39057] = 8'b1011000;
DRAM[39058] = 8'b1010101;
DRAM[39059] = 8'b1010101;
DRAM[39060] = 8'b1011000;
DRAM[39061] = 8'b1011100;
DRAM[39062] = 8'b1011111;
DRAM[39063] = 8'b1100000;
DRAM[39064] = 8'b1101011;
DRAM[39065] = 8'b1101100;
DRAM[39066] = 8'b1100101;
DRAM[39067] = 8'b1100101;
DRAM[39068] = 8'b1110101;
DRAM[39069] = 8'b10000101;
DRAM[39070] = 8'b10011000;
DRAM[39071] = 8'b10101111;
DRAM[39072] = 8'b1100110;
DRAM[39073] = 8'b1011001;
DRAM[39074] = 8'b10000001;
DRAM[39075] = 8'b10010101;
DRAM[39076] = 8'b10100010;
DRAM[39077] = 8'b11000001;
DRAM[39078] = 8'b11000110;
DRAM[39079] = 8'b11001001;
DRAM[39080] = 8'b11011101;
DRAM[39081] = 8'b11100001;
DRAM[39082] = 8'b11100111;
DRAM[39083] = 8'b11101101;
DRAM[39084] = 8'b11101111;
DRAM[39085] = 8'b11101111;
DRAM[39086] = 8'b11101111;
DRAM[39087] = 8'b11101110;
DRAM[39088] = 8'b11101000;
DRAM[39089] = 8'b11100100;
DRAM[39090] = 8'b11010101;
DRAM[39091] = 8'b11000010;
DRAM[39092] = 8'b11000000;
DRAM[39093] = 8'b11001000;
DRAM[39094] = 8'b11000010;
DRAM[39095] = 8'b10110011;
DRAM[39096] = 8'b10111010;
DRAM[39097] = 8'b10111010;
DRAM[39098] = 8'b10111100;
DRAM[39099] = 8'b11000000;
DRAM[39100] = 8'b11000010;
DRAM[39101] = 8'b10111110;
DRAM[39102] = 8'b10110100;
DRAM[39103] = 8'b10101100;
DRAM[39104] = 8'b10011101;
DRAM[39105] = 8'b10100110;
DRAM[39106] = 8'b10110100;
DRAM[39107] = 8'b11000101;
DRAM[39108] = 8'b11010110;
DRAM[39109] = 8'b11100011;
DRAM[39110] = 8'b11101000;
DRAM[39111] = 8'b11100111;
DRAM[39112] = 8'b11101011;
DRAM[39113] = 8'b11100101;
DRAM[39114] = 8'b11011101;
DRAM[39115] = 8'b11010011;
DRAM[39116] = 8'b11001001;
DRAM[39117] = 8'b10111101;
DRAM[39118] = 8'b10110001;
DRAM[39119] = 8'b10101001;
DRAM[39120] = 8'b10011001;
DRAM[39121] = 8'b10010011;
DRAM[39122] = 8'b10001100;
DRAM[39123] = 8'b10001011;
DRAM[39124] = 8'b10001101;
DRAM[39125] = 8'b10010000;
DRAM[39126] = 8'b10001110;
DRAM[39127] = 8'b10001100;
DRAM[39128] = 8'b10010001;
DRAM[39129] = 8'b10010000;
DRAM[39130] = 8'b10010000;
DRAM[39131] = 8'b10001111;
DRAM[39132] = 8'b10001110;
DRAM[39133] = 8'b10001100;
DRAM[39134] = 8'b10001011;
DRAM[39135] = 8'b10001010;
DRAM[39136] = 8'b10001001;
DRAM[39137] = 8'b10001001;
DRAM[39138] = 8'b10001001;
DRAM[39139] = 8'b10001000;
DRAM[39140] = 8'b10000111;
DRAM[39141] = 8'b10000110;
DRAM[39142] = 8'b10000100;
DRAM[39143] = 8'b10000011;
DRAM[39144] = 8'b10000001;
DRAM[39145] = 8'b10000000;
DRAM[39146] = 8'b1111111;
DRAM[39147] = 8'b1111110;
DRAM[39148] = 8'b1111110;
DRAM[39149] = 8'b1111110;
DRAM[39150] = 8'b1111110;
DRAM[39151] = 8'b1111111;
DRAM[39152] = 8'b1111101;
DRAM[39153] = 8'b1111101;
DRAM[39154] = 8'b1111101;
DRAM[39155] = 8'b1111110;
DRAM[39156] = 8'b1111110;
DRAM[39157] = 8'b1111111;
DRAM[39158] = 8'b1111111;
DRAM[39159] = 8'b1111111;
DRAM[39160] = 8'b10000000;
DRAM[39161] = 8'b10000000;
DRAM[39162] = 8'b1111111;
DRAM[39163] = 8'b1111110;
DRAM[39164] = 8'b1111110;
DRAM[39165] = 8'b1111101;
DRAM[39166] = 8'b1111100;
DRAM[39167] = 8'b1111100;
DRAM[39168] = 8'b10011010;
DRAM[39169] = 8'b10011010;
DRAM[39170] = 8'b10011010;
DRAM[39171] = 8'b10011011;
DRAM[39172] = 8'b10011011;
DRAM[39173] = 8'b10011011;
DRAM[39174] = 8'b10011100;
DRAM[39175] = 8'b10011100;
DRAM[39176] = 8'b10011101;
DRAM[39177] = 8'b10011101;
DRAM[39178] = 8'b10011101;
DRAM[39179] = 8'b10011101;
DRAM[39180] = 8'b10011110;
DRAM[39181] = 8'b10011111;
DRAM[39182] = 8'b10100000;
DRAM[39183] = 8'b10100001;
DRAM[39184] = 8'b10100001;
DRAM[39185] = 8'b10100001;
DRAM[39186] = 8'b10100010;
DRAM[39187] = 8'b10100010;
DRAM[39188] = 8'b10100011;
DRAM[39189] = 8'b10100100;
DRAM[39190] = 8'b10100101;
DRAM[39191] = 8'b10100101;
DRAM[39192] = 8'b10100101;
DRAM[39193] = 8'b10100100;
DRAM[39194] = 8'b10100100;
DRAM[39195] = 8'b10100100;
DRAM[39196] = 8'b10100100;
DRAM[39197] = 8'b10100101;
DRAM[39198] = 8'b10100110;
DRAM[39199] = 8'b10100111;
DRAM[39200] = 8'b10101000;
DRAM[39201] = 8'b10101000;
DRAM[39202] = 8'b10100111;
DRAM[39203] = 8'b10100110;
DRAM[39204] = 8'b10100110;
DRAM[39205] = 8'b10100101;
DRAM[39206] = 8'b10100100;
DRAM[39207] = 8'b10100100;
DRAM[39208] = 8'b10100100;
DRAM[39209] = 8'b10100010;
DRAM[39210] = 8'b10100001;
DRAM[39211] = 8'b10100100;
DRAM[39212] = 8'b10100101;
DRAM[39213] = 8'b10100100;
DRAM[39214] = 8'b10100111;
DRAM[39215] = 8'b10101100;
DRAM[39216] = 8'b10110011;
DRAM[39217] = 8'b11000111;
DRAM[39218] = 8'b11100010;
DRAM[39219] = 8'b11110100;
DRAM[39220] = 8'b11111010;
DRAM[39221] = 8'b11111011;
DRAM[39222] = 8'b11111100;
DRAM[39223] = 8'b11111110;
DRAM[39224] = 8'b11111101;
DRAM[39225] = 8'b11111100;
DRAM[39226] = 8'b11111101;
DRAM[39227] = 8'b11111101;
DRAM[39228] = 8'b11111110;
DRAM[39229] = 8'b11111100;
DRAM[39230] = 8'b11111000;
DRAM[39231] = 8'b11110100;
DRAM[39232] = 8'b11101000;
DRAM[39233] = 8'b11011110;
DRAM[39234] = 8'b11010001;
DRAM[39235] = 8'b11000111;
DRAM[39236] = 8'b11000010;
DRAM[39237] = 8'b10111101;
DRAM[39238] = 8'b10110110;
DRAM[39239] = 8'b10110000;
DRAM[39240] = 8'b10101011;
DRAM[39241] = 8'b10101110;
DRAM[39242] = 8'b10101110;
DRAM[39243] = 8'b10101100;
DRAM[39244] = 8'b10101110;
DRAM[39245] = 8'b10110011;
DRAM[39246] = 8'b10110011;
DRAM[39247] = 8'b10101110;
DRAM[39248] = 8'b10100101;
DRAM[39249] = 8'b10011101;
DRAM[39250] = 8'b10011000;
DRAM[39251] = 8'b10011101;
DRAM[39252] = 8'b10100011;
DRAM[39253] = 8'b10100101;
DRAM[39254] = 8'b10100101;
DRAM[39255] = 8'b10100111;
DRAM[39256] = 8'b10100110;
DRAM[39257] = 8'b10101011;
DRAM[39258] = 8'b10101100;
DRAM[39259] = 8'b10101001;
DRAM[39260] = 8'b10101100;
DRAM[39261] = 8'b10110110;
DRAM[39262] = 8'b10111111;
DRAM[39263] = 8'b11000010;
DRAM[39264] = 8'b11001000;
DRAM[39265] = 8'b11000011;
DRAM[39266] = 8'b10111110;
DRAM[39267] = 8'b10111011;
DRAM[39268] = 8'b10111010;
DRAM[39269] = 8'b10111011;
DRAM[39270] = 8'b10111100;
DRAM[39271] = 8'b10111011;
DRAM[39272] = 8'b10111001;
DRAM[39273] = 8'b10111110;
DRAM[39274] = 8'b10111010;
DRAM[39275] = 8'b10110010;
DRAM[39276] = 8'b10110101;
DRAM[39277] = 8'b11000000;
DRAM[39278] = 8'b10111111;
DRAM[39279] = 8'b10110100;
DRAM[39280] = 8'b10110011;
DRAM[39281] = 8'b10111100;
DRAM[39282] = 8'b11001011;
DRAM[39283] = 8'b11011010;
DRAM[39284] = 8'b11011110;
DRAM[39285] = 8'b11011101;
DRAM[39286] = 8'b11011110;
DRAM[39287] = 8'b11100010;
DRAM[39288] = 8'b11011011;
DRAM[39289] = 8'b11011100;
DRAM[39290] = 8'b11100101;
DRAM[39291] = 8'b11101010;
DRAM[39292] = 8'b11100110;
DRAM[39293] = 8'b11100100;
DRAM[39294] = 8'b11011010;
DRAM[39295] = 8'b11001001;
DRAM[39296] = 8'b10111111;
DRAM[39297] = 8'b11000011;
DRAM[39298] = 8'b10101111;
DRAM[39299] = 8'b10101101;
DRAM[39300] = 8'b10011101;
DRAM[39301] = 8'b1101100;
DRAM[39302] = 8'b1011010;
DRAM[39303] = 8'b1100000;
DRAM[39304] = 8'b10000111;
DRAM[39305] = 8'b10000010;
DRAM[39306] = 8'b1110111;
DRAM[39307] = 8'b1101000;
DRAM[39308] = 8'b1011010;
DRAM[39309] = 8'b1010001;
DRAM[39310] = 8'b1001101;
DRAM[39311] = 8'b1001011;
DRAM[39312] = 8'b1001100;
DRAM[39313] = 8'b1001001;
DRAM[39314] = 8'b1000110;
DRAM[39315] = 8'b1000110;
DRAM[39316] = 8'b1001001;
DRAM[39317] = 8'b1001100;
DRAM[39318] = 8'b1001110;
DRAM[39319] = 8'b1001111;
DRAM[39320] = 8'b1010000;
DRAM[39321] = 8'b1010011;
DRAM[39322] = 8'b1001101;
DRAM[39323] = 8'b1001110;
DRAM[39324] = 8'b1011110;
DRAM[39325] = 8'b1101111;
DRAM[39326] = 8'b10000110;
DRAM[39327] = 8'b10100001;
DRAM[39328] = 8'b1111111;
DRAM[39329] = 8'b1010101;
DRAM[39330] = 8'b1100100;
DRAM[39331] = 8'b1111110;
DRAM[39332] = 8'b10010111;
DRAM[39333] = 8'b10110110;
DRAM[39334] = 8'b11000000;
DRAM[39335] = 8'b11001110;
DRAM[39336] = 8'b11100010;
DRAM[39337] = 8'b11100011;
DRAM[39338] = 8'b11100101;
DRAM[39339] = 8'b11101001;
DRAM[39340] = 8'b11101101;
DRAM[39341] = 8'b11101110;
DRAM[39342] = 8'b11101101;
DRAM[39343] = 8'b11101100;
DRAM[39344] = 8'b11100100;
DRAM[39345] = 8'b11100100;
DRAM[39346] = 8'b11011100;
DRAM[39347] = 8'b11001110;
DRAM[39348] = 8'b11001000;
DRAM[39349] = 8'b11001001;
DRAM[39350] = 8'b11001000;
DRAM[39351] = 8'b11000001;
DRAM[39352] = 8'b10111101;
DRAM[39353] = 8'b10111001;
DRAM[39354] = 8'b10110101;
DRAM[39355] = 8'b10110110;
DRAM[39356] = 8'b10111000;
DRAM[39357] = 8'b10111000;
DRAM[39358] = 8'b10110100;
DRAM[39359] = 8'b10110000;
DRAM[39360] = 8'b10101111;
DRAM[39361] = 8'b10111000;
DRAM[39362] = 8'b11000100;
DRAM[39363] = 8'b11001110;
DRAM[39364] = 8'b11010101;
DRAM[39365] = 8'b11011011;
DRAM[39366] = 8'b11011111;
DRAM[39367] = 8'b11100010;
DRAM[39368] = 8'b11010101;
DRAM[39369] = 8'b11100100;
DRAM[39370] = 8'b11110011;
DRAM[39371] = 8'b11110010;
DRAM[39372] = 8'b11100011;
DRAM[39373] = 8'b11010000;
DRAM[39374] = 8'b11000101;
DRAM[39375] = 8'b11000011;
DRAM[39376] = 8'b10110010;
DRAM[39377] = 8'b10101011;
DRAM[39378] = 8'b10100010;
DRAM[39379] = 8'b10011101;
DRAM[39380] = 8'b10011011;
DRAM[39381] = 8'b10011010;
DRAM[39382] = 8'b10010110;
DRAM[39383] = 8'b10010010;
DRAM[39384] = 8'b10001101;
DRAM[39385] = 8'b10001100;
DRAM[39386] = 8'b10001010;
DRAM[39387] = 8'b10001001;
DRAM[39388] = 8'b10001001;
DRAM[39389] = 8'b10001011;
DRAM[39390] = 8'b10001100;
DRAM[39391] = 8'b10001101;
DRAM[39392] = 8'b10001001;
DRAM[39393] = 8'b10001001;
DRAM[39394] = 8'b10001001;
DRAM[39395] = 8'b10001000;
DRAM[39396] = 8'b10000111;
DRAM[39397] = 8'b10000101;
DRAM[39398] = 8'b10000100;
DRAM[39399] = 8'b10000011;
DRAM[39400] = 8'b10000001;
DRAM[39401] = 8'b10000000;
DRAM[39402] = 8'b1111111;
DRAM[39403] = 8'b1111110;
DRAM[39404] = 8'b1111110;
DRAM[39405] = 8'b1111110;
DRAM[39406] = 8'b1111110;
DRAM[39407] = 8'b1111111;
DRAM[39408] = 8'b1111101;
DRAM[39409] = 8'b1111101;
DRAM[39410] = 8'b1111110;
DRAM[39411] = 8'b1111110;
DRAM[39412] = 8'b1111110;
DRAM[39413] = 8'b1111111;
DRAM[39414] = 8'b1111111;
DRAM[39415] = 8'b1111111;
DRAM[39416] = 8'b10000000;
DRAM[39417] = 8'b10000000;
DRAM[39418] = 8'b1111111;
DRAM[39419] = 8'b1111111;
DRAM[39420] = 8'b1111110;
DRAM[39421] = 8'b1111101;
DRAM[39422] = 8'b1111100;
DRAM[39423] = 8'b1111100;
DRAM[39424] = 8'b10011010;
DRAM[39425] = 8'b10011010;
DRAM[39426] = 8'b10011010;
DRAM[39427] = 8'b10011010;
DRAM[39428] = 8'b10011011;
DRAM[39429] = 8'b10011011;
DRAM[39430] = 8'b10011011;
DRAM[39431] = 8'b10011100;
DRAM[39432] = 8'b10011110;
DRAM[39433] = 8'b10011110;
DRAM[39434] = 8'b10011101;
DRAM[39435] = 8'b10011101;
DRAM[39436] = 8'b10011101;
DRAM[39437] = 8'b10011110;
DRAM[39438] = 8'b10011111;
DRAM[39439] = 8'b10011111;
DRAM[39440] = 8'b10100001;
DRAM[39441] = 8'b10100001;
DRAM[39442] = 8'b10100001;
DRAM[39443] = 8'b10100010;
DRAM[39444] = 8'b10100011;
DRAM[39445] = 8'b10100100;
DRAM[39446] = 8'b10100100;
DRAM[39447] = 8'b10100101;
DRAM[39448] = 8'b10100101;
DRAM[39449] = 8'b10100100;
DRAM[39450] = 8'b10100100;
DRAM[39451] = 8'b10100100;
DRAM[39452] = 8'b10100100;
DRAM[39453] = 8'b10100101;
DRAM[39454] = 8'b10100110;
DRAM[39455] = 8'b10100111;
DRAM[39456] = 8'b10101000;
DRAM[39457] = 8'b10101000;
DRAM[39458] = 8'b10100111;
DRAM[39459] = 8'b10100110;
DRAM[39460] = 8'b10100110;
DRAM[39461] = 8'b10100101;
DRAM[39462] = 8'b10100100;
DRAM[39463] = 8'b10100100;
DRAM[39464] = 8'b10100101;
DRAM[39465] = 8'b10100011;
DRAM[39466] = 8'b10100100;
DRAM[39467] = 8'b10100110;
DRAM[39468] = 8'b10100110;
DRAM[39469] = 8'b10100110;
DRAM[39470] = 8'b10101010;
DRAM[39471] = 8'b10110001;
DRAM[39472] = 8'b10111100;
DRAM[39473] = 8'b11011001;
DRAM[39474] = 8'b11110101;
DRAM[39475] = 8'b11111100;
DRAM[39476] = 8'b11111001;
DRAM[39477] = 8'b11111010;
DRAM[39478] = 8'b11111101;
DRAM[39479] = 8'b11111100;
DRAM[39480] = 8'b11111101;
DRAM[39481] = 8'b11111101;
DRAM[39482] = 8'b11111101;
DRAM[39483] = 8'b11111110;
DRAM[39484] = 8'b11111110;
DRAM[39485] = 8'b11111100;
DRAM[39486] = 8'b11111000;
DRAM[39487] = 8'b11110101;
DRAM[39488] = 8'b11100110;
DRAM[39489] = 8'b11011111;
DRAM[39490] = 8'b11010101;
DRAM[39491] = 8'b11001011;
DRAM[39492] = 8'b11000100;
DRAM[39493] = 8'b10111110;
DRAM[39494] = 8'b10111001;
DRAM[39495] = 8'b10110110;
DRAM[39496] = 8'b10100111;
DRAM[39497] = 8'b10101000;
DRAM[39498] = 8'b10100110;
DRAM[39499] = 8'b10100100;
DRAM[39500] = 8'b10100110;
DRAM[39501] = 8'b10101011;
DRAM[39502] = 8'b10101100;
DRAM[39503] = 8'b10101001;
DRAM[39504] = 8'b10100011;
DRAM[39505] = 8'b10011101;
DRAM[39506] = 8'b10011101;
DRAM[39507] = 8'b10100100;
DRAM[39508] = 8'b10101001;
DRAM[39509] = 8'b10101000;
DRAM[39510] = 8'b10100100;
DRAM[39511] = 8'b10100010;
DRAM[39512] = 8'b10101001;
DRAM[39513] = 8'b10101001;
DRAM[39514] = 8'b10101001;
DRAM[39515] = 8'b10101101;
DRAM[39516] = 8'b10110111;
DRAM[39517] = 8'b11000010;
DRAM[39518] = 8'b11000110;
DRAM[39519] = 8'b11000100;
DRAM[39520] = 8'b11000111;
DRAM[39521] = 8'b11000100;
DRAM[39522] = 8'b11000001;
DRAM[39523] = 8'b11000010;
DRAM[39524] = 8'b11000101;
DRAM[39525] = 8'b11000101;
DRAM[39526] = 8'b11000000;
DRAM[39527] = 8'b10111011;
DRAM[39528] = 8'b10111001;
DRAM[39529] = 8'b11000010;
DRAM[39530] = 8'b10111100;
DRAM[39531] = 8'b10101100;
DRAM[39532] = 8'b10110000;
DRAM[39533] = 8'b11000011;
DRAM[39534] = 8'b11000011;
DRAM[39535] = 8'b10110011;
DRAM[39536] = 8'b10111100;
DRAM[39537] = 8'b11000111;
DRAM[39538] = 8'b11010011;
DRAM[39539] = 8'b11011011;
DRAM[39540] = 8'b11100001;
DRAM[39541] = 8'b11100011;
DRAM[39542] = 8'b11011110;
DRAM[39543] = 8'b11011000;
DRAM[39544] = 8'b11011001;
DRAM[39545] = 8'b11100010;
DRAM[39546] = 8'b11100001;
DRAM[39547] = 8'b11011111;
DRAM[39548] = 8'b11100001;
DRAM[39549] = 8'b11011000;
DRAM[39550] = 8'b11000110;
DRAM[39551] = 8'b10111011;
DRAM[39552] = 8'b10110101;
DRAM[39553] = 8'b10101110;
DRAM[39554] = 8'b10011100;
DRAM[39555] = 8'b10100001;
DRAM[39556] = 8'b10001000;
DRAM[39557] = 8'b1010001;
DRAM[39558] = 8'b1001110;
DRAM[39559] = 8'b1101001;
DRAM[39560] = 8'b10001011;
DRAM[39561] = 8'b1111011;
DRAM[39562] = 8'b1100101;
DRAM[39563] = 8'b1010100;
DRAM[39564] = 8'b1001010;
DRAM[39565] = 8'b1000101;
DRAM[39566] = 8'b1000010;
DRAM[39567] = 8'b1000000;
DRAM[39568] = 8'b111101;
DRAM[39569] = 8'b111010;
DRAM[39570] = 8'b110111;
DRAM[39571] = 8'b110111;
DRAM[39572] = 8'b111001;
DRAM[39573] = 8'b111100;
DRAM[39574] = 8'b111101;
DRAM[39575] = 8'b111101;
DRAM[39576] = 8'b110111;
DRAM[39577] = 8'b111011;
DRAM[39578] = 8'b110111;
DRAM[39579] = 8'b111001;
DRAM[39580] = 8'b1000110;
DRAM[39581] = 8'b1010111;
DRAM[39582] = 8'b1110010;
DRAM[39583] = 8'b10010011;
DRAM[39584] = 8'b10010010;
DRAM[39585] = 8'b1010010;
DRAM[39586] = 8'b1001000;
DRAM[39587] = 8'b1101010;
DRAM[39588] = 8'b10010001;
DRAM[39589] = 8'b10101101;
DRAM[39590] = 8'b10111011;
DRAM[39591] = 8'b11010000;
DRAM[39592] = 8'b11100011;
DRAM[39593] = 8'b11100010;
DRAM[39594] = 8'b11100010;
DRAM[39595] = 8'b11100100;
DRAM[39596] = 8'b11101001;
DRAM[39597] = 8'b11101101;
DRAM[39598] = 8'b11101111;
DRAM[39599] = 8'b11110000;
DRAM[39600] = 8'b11100100;
DRAM[39601] = 8'b11100110;
DRAM[39602] = 8'b11100100;
DRAM[39603] = 8'b11011011;
DRAM[39604] = 8'b11001111;
DRAM[39605] = 8'b11001000;
DRAM[39606] = 8'b11001000;
DRAM[39607] = 8'b11001011;
DRAM[39608] = 8'b10111111;
DRAM[39609] = 8'b10111010;
DRAM[39610] = 8'b10110101;
DRAM[39611] = 8'b10110100;
DRAM[39612] = 8'b10110111;
DRAM[39613] = 8'b10110111;
DRAM[39614] = 8'b10110100;
DRAM[39615] = 8'b10110000;
DRAM[39616] = 8'b10110011;
DRAM[39617] = 8'b10111101;
DRAM[39618] = 8'b11001010;
DRAM[39619] = 8'b11010010;
DRAM[39620] = 8'b11010101;
DRAM[39621] = 8'b11011000;
DRAM[39622] = 8'b11011111;
DRAM[39623] = 8'b11100110;
DRAM[39624] = 8'b11101001;
DRAM[39625] = 8'b11101100;
DRAM[39626] = 8'b11110000;
DRAM[39627] = 8'b11110000;
DRAM[39628] = 8'b11100110;
DRAM[39629] = 8'b11001110;
DRAM[39630] = 8'b10101111;
DRAM[39631] = 8'b10011001;
DRAM[39632] = 8'b10101100;
DRAM[39633] = 8'b10100111;
DRAM[39634] = 8'b10100001;
DRAM[39635] = 8'b10011110;
DRAM[39636] = 8'b10011111;
DRAM[39637] = 8'b10011111;
DRAM[39638] = 8'b10011101;
DRAM[39639] = 8'b10011010;
DRAM[39640] = 8'b10011100;
DRAM[39641] = 8'b10011000;
DRAM[39642] = 8'b10010011;
DRAM[39643] = 8'b10001111;
DRAM[39644] = 8'b10001011;
DRAM[39645] = 8'b10001011;
DRAM[39646] = 8'b10001011;
DRAM[39647] = 8'b10001100;
DRAM[39648] = 8'b10001010;
DRAM[39649] = 8'b10001001;
DRAM[39650] = 8'b10001000;
DRAM[39651] = 8'b10000111;
DRAM[39652] = 8'b10000110;
DRAM[39653] = 8'b10000101;
DRAM[39654] = 8'b10000100;
DRAM[39655] = 8'b10000011;
DRAM[39656] = 8'b10000001;
DRAM[39657] = 8'b10000000;
DRAM[39658] = 8'b1111111;
DRAM[39659] = 8'b1111110;
DRAM[39660] = 8'b1111110;
DRAM[39661] = 8'b1111110;
DRAM[39662] = 8'b1111110;
DRAM[39663] = 8'b1111111;
DRAM[39664] = 8'b1111101;
DRAM[39665] = 8'b1111110;
DRAM[39666] = 8'b1111110;
DRAM[39667] = 8'b1111110;
DRAM[39668] = 8'b1111111;
DRAM[39669] = 8'b1111111;
DRAM[39670] = 8'b1111111;
DRAM[39671] = 8'b1111111;
DRAM[39672] = 8'b10000000;
DRAM[39673] = 8'b10000000;
DRAM[39674] = 8'b10000000;
DRAM[39675] = 8'b1111111;
DRAM[39676] = 8'b1111110;
DRAM[39677] = 8'b1111101;
DRAM[39678] = 8'b1111101;
DRAM[39679] = 8'b1111100;
DRAM[39680] = 8'b10011001;
DRAM[39681] = 8'b10011001;
DRAM[39682] = 8'b10011010;
DRAM[39683] = 8'b10011010;
DRAM[39684] = 8'b10011010;
DRAM[39685] = 8'b10011011;
DRAM[39686] = 8'b10011011;
DRAM[39687] = 8'b10011011;
DRAM[39688] = 8'b10011111;
DRAM[39689] = 8'b10011111;
DRAM[39690] = 8'b10011110;
DRAM[39691] = 8'b10011101;
DRAM[39692] = 8'b10011101;
DRAM[39693] = 8'b10011101;
DRAM[39694] = 8'b10011110;
DRAM[39695] = 8'b10011110;
DRAM[39696] = 8'b10100000;
DRAM[39697] = 8'b10100000;
DRAM[39698] = 8'b10100001;
DRAM[39699] = 8'b10100010;
DRAM[39700] = 8'b10100011;
DRAM[39701] = 8'b10100011;
DRAM[39702] = 8'b10100100;
DRAM[39703] = 8'b10100100;
DRAM[39704] = 8'b10100101;
DRAM[39705] = 8'b10100100;
DRAM[39706] = 8'b10100100;
DRAM[39707] = 8'b10100100;
DRAM[39708] = 8'b10100100;
DRAM[39709] = 8'b10100101;
DRAM[39710] = 8'b10100110;
DRAM[39711] = 8'b10100111;
DRAM[39712] = 8'b10100111;
DRAM[39713] = 8'b10100111;
DRAM[39714] = 8'b10100111;
DRAM[39715] = 8'b10100110;
DRAM[39716] = 8'b10100110;
DRAM[39717] = 8'b10100101;
DRAM[39718] = 8'b10100101;
DRAM[39719] = 8'b10100101;
DRAM[39720] = 8'b10101001;
DRAM[39721] = 8'b10100111;
DRAM[39722] = 8'b10100110;
DRAM[39723] = 8'b10101000;
DRAM[39724] = 8'b10100111;
DRAM[39725] = 8'b10100110;
DRAM[39726] = 8'b10101100;
DRAM[39727] = 8'b10110100;
DRAM[39728] = 8'b11010000;
DRAM[39729] = 8'b11101100;
DRAM[39730] = 8'b11111111;
DRAM[39731] = 8'b11111110;
DRAM[39732] = 8'b11111001;
DRAM[39733] = 8'b11111101;
DRAM[39734] = 8'b11111111;
DRAM[39735] = 8'b11111011;
DRAM[39736] = 8'b11111110;
DRAM[39737] = 8'b11111101;
DRAM[39738] = 8'b11111101;
DRAM[39739] = 8'b11111110;
DRAM[39740] = 8'b11111110;
DRAM[39741] = 8'b11111100;
DRAM[39742] = 8'b11111000;
DRAM[39743] = 8'b11110101;
DRAM[39744] = 8'b11101000;
DRAM[39745] = 8'b11100011;
DRAM[39746] = 8'b11011010;
DRAM[39747] = 8'b11010000;
DRAM[39748] = 8'b11000110;
DRAM[39749] = 8'b10111111;
DRAM[39750] = 8'b10111011;
DRAM[39751] = 8'b10111001;
DRAM[39752] = 8'b10110010;
DRAM[39753] = 8'b10110000;
DRAM[39754] = 8'b10101100;
DRAM[39755] = 8'b10101001;
DRAM[39756] = 8'b10101010;
DRAM[39757] = 8'b10101101;
DRAM[39758] = 8'b10101110;
DRAM[39759] = 8'b10101101;
DRAM[39760] = 8'b10100110;
DRAM[39761] = 8'b10100101;
DRAM[39762] = 8'b10100110;
DRAM[39763] = 8'b10101010;
DRAM[39764] = 8'b10101001;
DRAM[39765] = 8'b10100101;
DRAM[39766] = 8'b10100011;
DRAM[39767] = 8'b10100101;
DRAM[39768] = 8'b10100000;
DRAM[39769] = 8'b10100001;
DRAM[39770] = 8'b10100101;
DRAM[39771] = 8'b10101100;
DRAM[39772] = 8'b10110100;
DRAM[39773] = 8'b10111001;
DRAM[39774] = 8'b10110111;
DRAM[39775] = 8'b10110010;
DRAM[39776] = 8'b11000010;
DRAM[39777] = 8'b11000011;
DRAM[39778] = 8'b11000101;
DRAM[39779] = 8'b11000111;
DRAM[39780] = 8'b11000111;
DRAM[39781] = 8'b11000100;
DRAM[39782] = 8'b10111110;
DRAM[39783] = 8'b10111001;
DRAM[39784] = 8'b10110101;
DRAM[39785] = 8'b11000001;
DRAM[39786] = 8'b11000001;
DRAM[39787] = 8'b10110100;
DRAM[39788] = 8'b10110000;
DRAM[39789] = 8'b10111011;
DRAM[39790] = 8'b11000100;
DRAM[39791] = 8'b11000101;
DRAM[39792] = 8'b11001011;
DRAM[39793] = 8'b11010100;
DRAM[39794] = 8'b11011001;
DRAM[39795] = 8'b11011010;
DRAM[39796] = 8'b11011110;
DRAM[39797] = 8'b11100010;
DRAM[39798] = 8'b11011011;
DRAM[39799] = 8'b11001110;
DRAM[39800] = 8'b11010100;
DRAM[39801] = 8'b11100001;
DRAM[39802] = 8'b11011011;
DRAM[39803] = 8'b11010100;
DRAM[39804] = 8'b11011100;
DRAM[39805] = 8'b11010001;
DRAM[39806] = 8'b10111010;
DRAM[39807] = 8'b10110111;
DRAM[39808] = 8'b10110000;
DRAM[39809] = 8'b10100100;
DRAM[39810] = 8'b10001111;
DRAM[39811] = 8'b10001001;
DRAM[39812] = 8'b1100110;
DRAM[39813] = 8'b111000;
DRAM[39814] = 8'b1001010;
DRAM[39815] = 8'b1101101;
DRAM[39816] = 8'b1111111;
DRAM[39817] = 8'b1101100;
DRAM[39818] = 8'b1010100;
DRAM[39819] = 8'b1000101;
DRAM[39820] = 8'b111101;
DRAM[39821] = 8'b110111;
DRAM[39822] = 8'b110100;
DRAM[39823] = 8'b110011;
DRAM[39824] = 8'b101100;
DRAM[39825] = 8'b101001;
DRAM[39826] = 8'b100110;
DRAM[39827] = 8'b100110;
DRAM[39828] = 8'b100111;
DRAM[39829] = 8'b101001;
DRAM[39830] = 8'b101001;
DRAM[39831] = 8'b101001;
DRAM[39832] = 8'b100100;
DRAM[39833] = 8'b101000;
DRAM[39834] = 8'b100101;
DRAM[39835] = 8'b100101;
DRAM[39836] = 8'b101111;
DRAM[39837] = 8'b111011;
DRAM[39838] = 8'b1011000;
DRAM[39839] = 8'b1111100;
DRAM[39840] = 8'b10001101;
DRAM[39841] = 8'b1011000;
DRAM[39842] = 8'b1000101;
DRAM[39843] = 8'b1100100;
DRAM[39844] = 8'b10001101;
DRAM[39845] = 8'b10100111;
DRAM[39846] = 8'b10110111;
DRAM[39847] = 8'b11001011;
DRAM[39848] = 8'b11011001;
DRAM[39849] = 8'b11011011;
DRAM[39850] = 8'b11011110;
DRAM[39851] = 8'b11011111;
DRAM[39852] = 8'b11100000;
DRAM[39853] = 8'b11100101;
DRAM[39854] = 8'b11101110;
DRAM[39855] = 8'b11110101;
DRAM[39856] = 8'b11101001;
DRAM[39857] = 8'b11101000;
DRAM[39858] = 8'b11100111;
DRAM[39859] = 8'b11100010;
DRAM[39860] = 8'b11010101;
DRAM[39861] = 8'b11001000;
DRAM[39862] = 8'b11000110;
DRAM[39863] = 8'b11001011;
DRAM[39864] = 8'b11000010;
DRAM[39865] = 8'b11000000;
DRAM[39866] = 8'b10111110;
DRAM[39867] = 8'b10111110;
DRAM[39868] = 8'b10111110;
DRAM[39869] = 8'b10111011;
DRAM[39870] = 8'b10110100;
DRAM[39871] = 8'b10101110;
DRAM[39872] = 8'b10111000;
DRAM[39873] = 8'b10111110;
DRAM[39874] = 8'b11001001;
DRAM[39875] = 8'b11010100;
DRAM[39876] = 8'b11011001;
DRAM[39877] = 8'b11011100;
DRAM[39878] = 8'b11100011;
DRAM[39879] = 8'b11101010;
DRAM[39880] = 8'b11100110;
DRAM[39881] = 8'b11011110;
DRAM[39882] = 8'b11010111;
DRAM[39883] = 8'b11011010;
DRAM[39884] = 8'b11011100;
DRAM[39885] = 8'b11001111;
DRAM[39886] = 8'b10110100;
DRAM[39887] = 8'b10011100;
DRAM[39888] = 8'b10011010;
DRAM[39889] = 8'b10010111;
DRAM[39890] = 8'b10010100;
DRAM[39891] = 8'b10010100;
DRAM[39892] = 8'b10010110;
DRAM[39893] = 8'b10011001;
DRAM[39894] = 8'b10011001;
DRAM[39895] = 8'b10011000;
DRAM[39896] = 8'b10100001;
DRAM[39897] = 8'b10011111;
DRAM[39898] = 8'b10011010;
DRAM[39899] = 8'b10010101;
DRAM[39900] = 8'b10010001;
DRAM[39901] = 8'b10001110;
DRAM[39902] = 8'b10001101;
DRAM[39903] = 8'b10001100;
DRAM[39904] = 8'b10001010;
DRAM[39905] = 8'b10001001;
DRAM[39906] = 8'b10001000;
DRAM[39907] = 8'b10000110;
DRAM[39908] = 8'b10000101;
DRAM[39909] = 8'b10000100;
DRAM[39910] = 8'b10000100;
DRAM[39911] = 8'b10000100;
DRAM[39912] = 8'b10000001;
DRAM[39913] = 8'b10000000;
DRAM[39914] = 8'b1111111;
DRAM[39915] = 8'b1111110;
DRAM[39916] = 8'b1111110;
DRAM[39917] = 8'b1111110;
DRAM[39918] = 8'b1111110;
DRAM[39919] = 8'b1111111;
DRAM[39920] = 8'b1111110;
DRAM[39921] = 8'b1111110;
DRAM[39922] = 8'b1111110;
DRAM[39923] = 8'b1111111;
DRAM[39924] = 8'b1111111;
DRAM[39925] = 8'b1111111;
DRAM[39926] = 8'b10000000;
DRAM[39927] = 8'b10000000;
DRAM[39928] = 8'b10000001;
DRAM[39929] = 8'b10000001;
DRAM[39930] = 8'b10000000;
DRAM[39931] = 8'b1111111;
DRAM[39932] = 8'b1111110;
DRAM[39933] = 8'b1111110;
DRAM[39934] = 8'b1111101;
DRAM[39935] = 8'b1111101;
DRAM[39936] = 8'b10011001;
DRAM[39937] = 8'b10011001;
DRAM[39938] = 8'b10011001;
DRAM[39939] = 8'b10011010;
DRAM[39940] = 8'b10011010;
DRAM[39941] = 8'b10011010;
DRAM[39942] = 8'b10011011;
DRAM[39943] = 8'b10011011;
DRAM[39944] = 8'b10011111;
DRAM[39945] = 8'b10011111;
DRAM[39946] = 8'b10011110;
DRAM[39947] = 8'b10011101;
DRAM[39948] = 8'b10011101;
DRAM[39949] = 8'b10011101;
DRAM[39950] = 8'b10011110;
DRAM[39951] = 8'b10011110;
DRAM[39952] = 8'b10100000;
DRAM[39953] = 8'b10100000;
DRAM[39954] = 8'b10100001;
DRAM[39955] = 8'b10100001;
DRAM[39956] = 8'b10100010;
DRAM[39957] = 8'b10100011;
DRAM[39958] = 8'b10100100;
DRAM[39959] = 8'b10100100;
DRAM[39960] = 8'b10100101;
DRAM[39961] = 8'b10100100;
DRAM[39962] = 8'b10100100;
DRAM[39963] = 8'b10100100;
DRAM[39964] = 8'b10100100;
DRAM[39965] = 8'b10100101;
DRAM[39966] = 8'b10100110;
DRAM[39967] = 8'b10100111;
DRAM[39968] = 8'b10100111;
DRAM[39969] = 8'b10100111;
DRAM[39970] = 8'b10100110;
DRAM[39971] = 8'b10100110;
DRAM[39972] = 8'b10100110;
DRAM[39973] = 8'b10100110;
DRAM[39974] = 8'b10100101;
DRAM[39975] = 8'b10100101;
DRAM[39976] = 8'b10101001;
DRAM[39977] = 8'b10100111;
DRAM[39978] = 8'b10100110;
DRAM[39979] = 8'b10100110;
DRAM[39980] = 8'b10100100;
DRAM[39981] = 8'b10100101;
DRAM[39982] = 8'b10101111;
DRAM[39983] = 8'b10111001;
DRAM[39984] = 8'b11100110;
DRAM[39985] = 8'b11111000;
DRAM[39986] = 8'b11111111;
DRAM[39987] = 8'b11111100;
DRAM[39988] = 8'b11111001;
DRAM[39989] = 8'b11111111;
DRAM[39990] = 8'b11111111;
DRAM[39991] = 8'b11111010;
DRAM[39992] = 8'b11111110;
DRAM[39993] = 8'b11111110;
DRAM[39994] = 8'b11111110;
DRAM[39995] = 8'b11111111;
DRAM[39996] = 8'b11111111;
DRAM[39997] = 8'b11111101;
DRAM[39998] = 8'b11111001;
DRAM[39999] = 8'b11110101;
DRAM[40000] = 8'b11101101;
DRAM[40001] = 8'b11100111;
DRAM[40002] = 8'b11011110;
DRAM[40003] = 8'b11010011;
DRAM[40004] = 8'b11001001;
DRAM[40005] = 8'b11000001;
DRAM[40006] = 8'b10111011;
DRAM[40007] = 8'b10111000;
DRAM[40008] = 8'b10110111;
DRAM[40009] = 8'b10110001;
DRAM[40010] = 8'b10101011;
DRAM[40011] = 8'b10101000;
DRAM[40012] = 8'b10100111;
DRAM[40013] = 8'b10100110;
DRAM[40014] = 8'b10100110;
DRAM[40015] = 8'b10100111;
DRAM[40016] = 8'b10101111;
DRAM[40017] = 8'b10110000;
DRAM[40018] = 8'b10110010;
DRAM[40019] = 8'b10110000;
DRAM[40020] = 8'b10101001;
DRAM[40021] = 8'b10100011;
DRAM[40022] = 8'b10101000;
DRAM[40023] = 8'b10110001;
DRAM[40024] = 8'b10101001;
DRAM[40025] = 8'b10101010;
DRAM[40026] = 8'b10101100;
DRAM[40027] = 8'b10101110;
DRAM[40028] = 8'b10101111;
DRAM[40029] = 8'b10101110;
DRAM[40030] = 8'b10101110;
DRAM[40031] = 8'b10101111;
DRAM[40032] = 8'b10111000;
DRAM[40033] = 8'b10111111;
DRAM[40034] = 8'b11000101;
DRAM[40035] = 8'b11000101;
DRAM[40036] = 8'b10111110;
DRAM[40037] = 8'b10111000;
DRAM[40038] = 8'b10110101;
DRAM[40039] = 8'b10110101;
DRAM[40040] = 8'b10110110;
DRAM[40041] = 8'b10110110;
DRAM[40042] = 8'b10111000;
DRAM[40043] = 8'b10111010;
DRAM[40044] = 8'b10111001;
DRAM[40045] = 8'b10111011;
DRAM[40046] = 8'b11000101;
DRAM[40047] = 8'b11010001;
DRAM[40048] = 8'b11010011;
DRAM[40049] = 8'b11011001;
DRAM[40050] = 8'b11011001;
DRAM[40051] = 8'b11010110;
DRAM[40052] = 8'b11011001;
DRAM[40053] = 8'b11011111;
DRAM[40054] = 8'b11011001;
DRAM[40055] = 8'b11001101;
DRAM[40056] = 8'b11001110;
DRAM[40057] = 8'b11011011;
DRAM[40058] = 8'b11010100;
DRAM[40059] = 8'b11001111;
DRAM[40060] = 8'b11011010;
DRAM[40061] = 8'b11010011;
DRAM[40062] = 8'b11000000;
DRAM[40063] = 8'b10111111;
DRAM[40064] = 8'b10110011;
DRAM[40065] = 8'b10101010;
DRAM[40066] = 8'b10001111;
DRAM[40067] = 8'b1110101;
DRAM[40068] = 8'b1001001;
DRAM[40069] = 8'b101111;
DRAM[40070] = 8'b1010001;
DRAM[40071] = 8'b1101110;
DRAM[40072] = 8'b1110001;
DRAM[40073] = 8'b1011101;
DRAM[40074] = 8'b1000111;
DRAM[40075] = 8'b111000;
DRAM[40076] = 8'b101011;
DRAM[40077] = 8'b11111;
DRAM[40078] = 8'b11000;
DRAM[40079] = 8'b10111;
DRAM[40080] = 8'b10101;
DRAM[40081] = 8'b10011;
DRAM[40082] = 8'b10000;
DRAM[40083] = 8'b10000;
DRAM[40084] = 8'b10001;
DRAM[40085] = 8'b10010;
DRAM[40086] = 8'b10010;
DRAM[40087] = 8'b10001;
DRAM[40088] = 8'b1111;
DRAM[40089] = 8'b10011;
DRAM[40090] = 8'b10000;
DRAM[40091] = 8'b1111;
DRAM[40092] = 8'b10100;
DRAM[40093] = 8'b11010;
DRAM[40094] = 8'b110011;
DRAM[40095] = 8'b1011000;
DRAM[40096] = 8'b1111111;
DRAM[40097] = 8'b1101001;
DRAM[40098] = 8'b1010011;
DRAM[40099] = 8'b1100001;
DRAM[40100] = 8'b10000001;
DRAM[40101] = 8'b10011011;
DRAM[40102] = 8'b10110010;
DRAM[40103] = 8'b10111111;
DRAM[40104] = 8'b11001010;
DRAM[40105] = 8'b11010010;
DRAM[40106] = 8'b11011000;
DRAM[40107] = 8'b11010111;
DRAM[40108] = 8'b11010011;
DRAM[40109] = 8'b11010110;
DRAM[40110] = 8'b11100100;
DRAM[40111] = 8'b11110001;
DRAM[40112] = 8'b11101110;
DRAM[40113] = 8'b11101001;
DRAM[40114] = 8'b11100101;
DRAM[40115] = 8'b11100010;
DRAM[40116] = 8'b11011011;
DRAM[40117] = 8'b11001111;
DRAM[40118] = 8'b11001010;
DRAM[40119] = 8'b11001011;
DRAM[40120] = 8'b11001001;
DRAM[40121] = 8'b11001001;
DRAM[40122] = 8'b11000110;
DRAM[40123] = 8'b11000011;
DRAM[40124] = 8'b10111110;
DRAM[40125] = 8'b10111001;
DRAM[40126] = 8'b10110100;
DRAM[40127] = 8'b10110010;
DRAM[40128] = 8'b11000100;
DRAM[40129] = 8'b11000100;
DRAM[40130] = 8'b11001010;
DRAM[40131] = 8'b11010101;
DRAM[40132] = 8'b11011101;
DRAM[40133] = 8'b11011110;
DRAM[40134] = 8'b11100000;
DRAM[40135] = 8'b11100100;
DRAM[40136] = 8'b11011101;
DRAM[40137] = 8'b11011110;
DRAM[40138] = 8'b11011101;
DRAM[40139] = 8'b11011001;
DRAM[40140] = 8'b11010010;
DRAM[40141] = 8'b11001001;
DRAM[40142] = 8'b11000010;
DRAM[40143] = 8'b10111101;
DRAM[40144] = 8'b10011101;
DRAM[40145] = 8'b10011010;
DRAM[40146] = 8'b10010111;
DRAM[40147] = 8'b10010100;
DRAM[40148] = 8'b10010010;
DRAM[40149] = 8'b10010001;
DRAM[40150] = 8'b10010000;
DRAM[40151] = 8'b10001111;
DRAM[40152] = 8'b10001111;
DRAM[40153] = 8'b10010000;
DRAM[40154] = 8'b10010001;
DRAM[40155] = 8'b10010010;
DRAM[40156] = 8'b10010010;
DRAM[40157] = 8'b10010000;
DRAM[40158] = 8'b10001111;
DRAM[40159] = 8'b10001101;
DRAM[40160] = 8'b10001010;
DRAM[40161] = 8'b10001001;
DRAM[40162] = 8'b10000111;
DRAM[40163] = 8'b10000101;
DRAM[40164] = 8'b10000100;
DRAM[40165] = 8'b10000100;
DRAM[40166] = 8'b10000100;
DRAM[40167] = 8'b10000100;
DRAM[40168] = 8'b10000001;
DRAM[40169] = 8'b10000000;
DRAM[40170] = 8'b1111111;
DRAM[40171] = 8'b1111110;
DRAM[40172] = 8'b1111110;
DRAM[40173] = 8'b1111110;
DRAM[40174] = 8'b1111110;
DRAM[40175] = 8'b1111111;
DRAM[40176] = 8'b1111110;
DRAM[40177] = 8'b1111110;
DRAM[40178] = 8'b1111111;
DRAM[40179] = 8'b1111111;
DRAM[40180] = 8'b1111111;
DRAM[40181] = 8'b10000000;
DRAM[40182] = 8'b10000000;
DRAM[40183] = 8'b10000000;
DRAM[40184] = 8'b10000001;
DRAM[40185] = 8'b10000001;
DRAM[40186] = 8'b10000000;
DRAM[40187] = 8'b10000000;
DRAM[40188] = 8'b1111111;
DRAM[40189] = 8'b1111110;
DRAM[40190] = 8'b1111101;
DRAM[40191] = 8'b1111101;
DRAM[40192] = 8'b10011000;
DRAM[40193] = 8'b10011001;
DRAM[40194] = 8'b10011001;
DRAM[40195] = 8'b10011001;
DRAM[40196] = 8'b10011010;
DRAM[40197] = 8'b10011010;
DRAM[40198] = 8'b10011010;
DRAM[40199] = 8'b10011010;
DRAM[40200] = 8'b10011110;
DRAM[40201] = 8'b10011110;
DRAM[40202] = 8'b10011101;
DRAM[40203] = 8'b10011101;
DRAM[40204] = 8'b10011101;
DRAM[40205] = 8'b10011110;
DRAM[40206] = 8'b10011111;
DRAM[40207] = 8'b10011111;
DRAM[40208] = 8'b10011111;
DRAM[40209] = 8'b10100000;
DRAM[40210] = 8'b10100000;
DRAM[40211] = 8'b10100001;
DRAM[40212] = 8'b10100010;
DRAM[40213] = 8'b10100011;
DRAM[40214] = 8'b10100011;
DRAM[40215] = 8'b10100011;
DRAM[40216] = 8'b10100101;
DRAM[40217] = 8'b10100100;
DRAM[40218] = 8'b10100100;
DRAM[40219] = 8'b10100100;
DRAM[40220] = 8'b10100100;
DRAM[40221] = 8'b10100101;
DRAM[40222] = 8'b10100110;
DRAM[40223] = 8'b10100111;
DRAM[40224] = 8'b10100110;
DRAM[40225] = 8'b10100110;
DRAM[40226] = 8'b10100110;
DRAM[40227] = 8'b10100110;
DRAM[40228] = 8'b10100110;
DRAM[40229] = 8'b10100110;
DRAM[40230] = 8'b10100110;
DRAM[40231] = 8'b10100110;
DRAM[40232] = 8'b10100110;
DRAM[40233] = 8'b10100100;
DRAM[40234] = 8'b10100100;
DRAM[40235] = 8'b10100100;
DRAM[40236] = 8'b10100101;
DRAM[40237] = 8'b10101011;
DRAM[40238] = 8'b10111010;
DRAM[40239] = 8'b11001001;
DRAM[40240] = 8'b11110110;
DRAM[40241] = 8'b11111101;
DRAM[40242] = 8'b11111111;
DRAM[40243] = 8'b11111011;
DRAM[40244] = 8'b11111011;
DRAM[40245] = 8'b11111111;
DRAM[40246] = 8'b11111111;
DRAM[40247] = 8'b11111011;
DRAM[40248] = 8'b11111110;
DRAM[40249] = 8'b11111110;
DRAM[40250] = 8'b11111110;
DRAM[40251] = 8'b11111111;
DRAM[40252] = 8'b11111111;
DRAM[40253] = 8'b11111101;
DRAM[40254] = 8'b11111001;
DRAM[40255] = 8'b11110110;
DRAM[40256] = 8'b11110000;
DRAM[40257] = 8'b11101001;
DRAM[40258] = 8'b11011111;
DRAM[40259] = 8'b11010101;
DRAM[40260] = 8'b11001100;
DRAM[40261] = 8'b11000100;
DRAM[40262] = 8'b10111100;
DRAM[40263] = 8'b10110111;
DRAM[40264] = 8'b10110011;
DRAM[40265] = 8'b10101100;
DRAM[40266] = 8'b10100101;
DRAM[40267] = 8'b10100010;
DRAM[40268] = 8'b10100000;
DRAM[40269] = 8'b10011100;
DRAM[40270] = 8'b10011011;
DRAM[40271] = 8'b10011100;
DRAM[40272] = 8'b10101101;
DRAM[40273] = 8'b10101110;
DRAM[40274] = 8'b10110000;
DRAM[40275] = 8'b10101110;
DRAM[40276] = 8'b10100110;
DRAM[40277] = 8'b10100000;
DRAM[40278] = 8'b10100110;
DRAM[40279] = 8'b10110001;
DRAM[40280] = 8'b10111000;
DRAM[40281] = 8'b10110110;
DRAM[40282] = 8'b10110100;
DRAM[40283] = 8'b10110001;
DRAM[40284] = 8'b10101100;
DRAM[40285] = 8'b10101011;
DRAM[40286] = 8'b10110010;
DRAM[40287] = 8'b10111011;
DRAM[40288] = 8'b10110011;
DRAM[40289] = 8'b10111011;
DRAM[40290] = 8'b11000001;
DRAM[40291] = 8'b10111110;
DRAM[40292] = 8'b10110101;
DRAM[40293] = 8'b10101110;
DRAM[40294] = 8'b10101111;
DRAM[40295] = 8'b10110011;
DRAM[40296] = 8'b11000001;
DRAM[40297] = 8'b10110011;
DRAM[40298] = 8'b10110000;
DRAM[40299] = 8'b11000000;
DRAM[40300] = 8'b11001101;
DRAM[40301] = 8'b11001110;
DRAM[40302] = 8'b11010000;
DRAM[40303] = 8'b11010101;
DRAM[40304] = 8'b11010011;
DRAM[40305] = 8'b11010101;
DRAM[40306] = 8'b11010101;
DRAM[40307] = 8'b11010101;
DRAM[40308] = 8'b11011000;
DRAM[40309] = 8'b11011100;
DRAM[40310] = 8'b11011010;
DRAM[40311] = 8'b11010100;
DRAM[40312] = 8'b11010111;
DRAM[40313] = 8'b11011011;
DRAM[40314] = 8'b11010101;
DRAM[40315] = 8'b11001111;
DRAM[40316] = 8'b11010010;
DRAM[40317] = 8'b11001110;
DRAM[40318] = 8'b11000010;
DRAM[40319] = 8'b10111100;
DRAM[40320] = 8'b10111001;
DRAM[40321] = 8'b10110011;
DRAM[40322] = 8'b10010110;
DRAM[40323] = 8'b1110001;
DRAM[40324] = 8'b1000000;
DRAM[40325] = 8'b110100;
DRAM[40326] = 8'b1011011;
DRAM[40327] = 8'b1101100;
DRAM[40328] = 8'b1011000;
DRAM[40329] = 8'b1000011;
DRAM[40330] = 8'b101110;
DRAM[40331] = 8'b100011;
DRAM[40332] = 8'b11001;
DRAM[40333] = 8'b1101;
DRAM[40334] = 8'b101;
DRAM[40335] = 8'b101;
DRAM[40336] = 8'b111;
DRAM[40337] = 8'b101;
DRAM[40338] = 8'b11;
DRAM[40339] = 8'b11;
DRAM[40340] = 8'b101;
DRAM[40341] = 8'b101;
DRAM[40342] = 8'b101;
DRAM[40343] = 8'b100;
DRAM[40344] = 8'b11;
DRAM[40345] = 8'b101;
DRAM[40346] = 8'b10;
DRAM[40347] = 8'b11;
DRAM[40348] = 8'b110;
DRAM[40349] = 8'b101;
DRAM[40350] = 8'b11001;
DRAM[40351] = 8'b111100;
DRAM[40352] = 8'b1110001;
DRAM[40353] = 8'b1110101;
DRAM[40354] = 8'b1011100;
DRAM[40355] = 8'b1011011;
DRAM[40356] = 8'b1110101;
DRAM[40357] = 8'b10001111;
DRAM[40358] = 8'b10101011;
DRAM[40359] = 8'b10110100;
DRAM[40360] = 8'b10111111;
DRAM[40361] = 8'b11001000;
DRAM[40362] = 8'b11010000;
DRAM[40363] = 8'b11001111;
DRAM[40364] = 8'b11001010;
DRAM[40365] = 8'b11001101;
DRAM[40366] = 8'b11011011;
DRAM[40367] = 8'b11101000;
DRAM[40368] = 8'b11101111;
DRAM[40369] = 8'b11101010;
DRAM[40370] = 8'b11100011;
DRAM[40371] = 8'b11011111;
DRAM[40372] = 8'b11011100;
DRAM[40373] = 8'b11011001;
DRAM[40374] = 8'b11010101;
DRAM[40375] = 8'b11010000;
DRAM[40376] = 8'b11010001;
DRAM[40377] = 8'b11001111;
DRAM[40378] = 8'b11001001;
DRAM[40379] = 8'b10111111;
DRAM[40380] = 8'b10110100;
DRAM[40381] = 8'b10110001;
DRAM[40382] = 8'b10110110;
DRAM[40383] = 8'b10111101;
DRAM[40384] = 8'b10111111;
DRAM[40385] = 8'b10111100;
DRAM[40386] = 8'b11000001;
DRAM[40387] = 8'b11010000;
DRAM[40388] = 8'b11011001;
DRAM[40389] = 8'b11011000;
DRAM[40390] = 8'b11011000;
DRAM[40391] = 8'b11011011;
DRAM[40392] = 8'b11100010;
DRAM[40393] = 8'b11011011;
DRAM[40394] = 8'b11010011;
DRAM[40395] = 8'b11001011;
DRAM[40396] = 8'b11000101;
DRAM[40397] = 8'b10111011;
DRAM[40398] = 8'b10101110;
DRAM[40399] = 8'b10100101;
DRAM[40400] = 8'b10100000;
DRAM[40401] = 8'b10011110;
DRAM[40402] = 8'b10011011;
DRAM[40403] = 8'b10011000;
DRAM[40404] = 8'b10010100;
DRAM[40405] = 8'b10010010;
DRAM[40406] = 8'b10010000;
DRAM[40407] = 8'b10001111;
DRAM[40408] = 8'b10001100;
DRAM[40409] = 8'b10001101;
DRAM[40410] = 8'b10010000;
DRAM[40411] = 8'b10010001;
DRAM[40412] = 8'b10010000;
DRAM[40413] = 8'b10001110;
DRAM[40414] = 8'b10001010;
DRAM[40415] = 8'b10001000;
DRAM[40416] = 8'b10001010;
DRAM[40417] = 8'b10001001;
DRAM[40418] = 8'b10000110;
DRAM[40419] = 8'b10000100;
DRAM[40420] = 8'b10000011;
DRAM[40421] = 8'b10000011;
DRAM[40422] = 8'b10000011;
DRAM[40423] = 8'b10000100;
DRAM[40424] = 8'b10000001;
DRAM[40425] = 8'b10000000;
DRAM[40426] = 8'b1111111;
DRAM[40427] = 8'b1111110;
DRAM[40428] = 8'b1111110;
DRAM[40429] = 8'b1111110;
DRAM[40430] = 8'b1111110;
DRAM[40431] = 8'b1111111;
DRAM[40432] = 8'b1111111;
DRAM[40433] = 8'b1111111;
DRAM[40434] = 8'b1111111;
DRAM[40435] = 8'b1111111;
DRAM[40436] = 8'b10000000;
DRAM[40437] = 8'b10000000;
DRAM[40438] = 8'b10000000;
DRAM[40439] = 8'b10000001;
DRAM[40440] = 8'b10000010;
DRAM[40441] = 8'b10000001;
DRAM[40442] = 8'b10000001;
DRAM[40443] = 8'b10000000;
DRAM[40444] = 8'b1111111;
DRAM[40445] = 8'b1111110;
DRAM[40446] = 8'b1111110;
DRAM[40447] = 8'b1111110;
DRAM[40448] = 8'b10011000;
DRAM[40449] = 8'b10011000;
DRAM[40450] = 8'b10011001;
DRAM[40451] = 8'b10011001;
DRAM[40452] = 8'b10011001;
DRAM[40453] = 8'b10011010;
DRAM[40454] = 8'b10011010;
DRAM[40455] = 8'b10011010;
DRAM[40456] = 8'b10011101;
DRAM[40457] = 8'b10011101;
DRAM[40458] = 8'b10011101;
DRAM[40459] = 8'b10011101;
DRAM[40460] = 8'b10011110;
DRAM[40461] = 8'b10011111;
DRAM[40462] = 8'b10100000;
DRAM[40463] = 8'b10100001;
DRAM[40464] = 8'b10011111;
DRAM[40465] = 8'b10011111;
DRAM[40466] = 8'b10100000;
DRAM[40467] = 8'b10100001;
DRAM[40468] = 8'b10100010;
DRAM[40469] = 8'b10100010;
DRAM[40470] = 8'b10100011;
DRAM[40471] = 8'b10100011;
DRAM[40472] = 8'b10100101;
DRAM[40473] = 8'b10100100;
DRAM[40474] = 8'b10100100;
DRAM[40475] = 8'b10100100;
DRAM[40476] = 8'b10100100;
DRAM[40477] = 8'b10100101;
DRAM[40478] = 8'b10100110;
DRAM[40479] = 8'b10100111;
DRAM[40480] = 8'b10100110;
DRAM[40481] = 8'b10100110;
DRAM[40482] = 8'b10100110;
DRAM[40483] = 8'b10100110;
DRAM[40484] = 8'b10100110;
DRAM[40485] = 8'b10100110;
DRAM[40486] = 8'b10100110;
DRAM[40487] = 8'b10100110;
DRAM[40488] = 8'b10100100;
DRAM[40489] = 8'b10100011;
DRAM[40490] = 8'b10100101;
DRAM[40491] = 8'b10101001;
DRAM[40492] = 8'b10101111;
DRAM[40493] = 8'b10111011;
DRAM[40494] = 8'b11010010;
DRAM[40495] = 8'b11100101;
DRAM[40496] = 8'b11111011;
DRAM[40497] = 8'b11111100;
DRAM[40498] = 8'b11111110;
DRAM[40499] = 8'b11111110;
DRAM[40500] = 8'b11111110;
DRAM[40501] = 8'b11111110;
DRAM[40502] = 8'b11111101;
DRAM[40503] = 8'b11111101;
DRAM[40504] = 8'b11111111;
DRAM[40505] = 8'b11111110;
DRAM[40506] = 8'b11111110;
DRAM[40507] = 8'b11111111;
DRAM[40508] = 8'b11111111;
DRAM[40509] = 8'b11111110;
DRAM[40510] = 8'b11111001;
DRAM[40511] = 8'b11110110;
DRAM[40512] = 8'b11110001;
DRAM[40513] = 8'b11101000;
DRAM[40514] = 8'b11011101;
DRAM[40515] = 8'b11010101;
DRAM[40516] = 8'b11001111;
DRAM[40517] = 8'b11001000;
DRAM[40518] = 8'b10111111;
DRAM[40519] = 8'b10110111;
DRAM[40520] = 8'b10111011;
DRAM[40521] = 8'b10110010;
DRAM[40522] = 8'b10101100;
DRAM[40523] = 8'b10101100;
DRAM[40524] = 8'b10101001;
DRAM[40525] = 8'b10100011;
DRAM[40526] = 8'b10100001;
DRAM[40527] = 8'b10100011;
DRAM[40528] = 8'b10100001;
DRAM[40529] = 8'b10100010;
DRAM[40530] = 8'b10100110;
DRAM[40531] = 8'b10101010;
DRAM[40532] = 8'b10101001;
DRAM[40533] = 8'b10100011;
DRAM[40534] = 8'b10100010;
DRAM[40535] = 8'b10100101;
DRAM[40536] = 8'b10101010;
DRAM[40537] = 8'b10101001;
DRAM[40538] = 8'b10101001;
DRAM[40539] = 8'b10101011;
DRAM[40540] = 8'b10101000;
DRAM[40541] = 8'b10100101;
DRAM[40542] = 8'b10101011;
DRAM[40543] = 8'b10110101;
DRAM[40544] = 8'b10111001;
DRAM[40545] = 8'b10111101;
DRAM[40546] = 8'b10111110;
DRAM[40547] = 8'b10111011;
DRAM[40548] = 8'b10110101;
DRAM[40549] = 8'b10110010;
DRAM[40550] = 8'b10110101;
DRAM[40551] = 8'b10111010;
DRAM[40552] = 8'b11000000;
DRAM[40553] = 8'b10111010;
DRAM[40554] = 8'b10111010;
DRAM[40555] = 8'b11000111;
DRAM[40556] = 8'b11010110;
DRAM[40557] = 8'b11011101;
DRAM[40558] = 8'b11011011;
DRAM[40559] = 8'b11011001;
DRAM[40560] = 8'b11010010;
DRAM[40561] = 8'b11010001;
DRAM[40562] = 8'b11010011;
DRAM[40563] = 8'b11011001;
DRAM[40564] = 8'b11011100;
DRAM[40565] = 8'b11011001;
DRAM[40566] = 8'b11010111;
DRAM[40567] = 8'b11011000;
DRAM[40568] = 8'b11011000;
DRAM[40569] = 8'b11010010;
DRAM[40570] = 8'b11010000;
DRAM[40571] = 8'b11001011;
DRAM[40572] = 8'b11000100;
DRAM[40573] = 8'b11000101;
DRAM[40574] = 8'b11000010;
DRAM[40575] = 8'b10110101;
DRAM[40576] = 8'b10111010;
DRAM[40577] = 8'b10110001;
DRAM[40578] = 8'b10011001;
DRAM[40579] = 8'b1111010;
DRAM[40580] = 8'b1001001;
DRAM[40581] = 8'b111010;
DRAM[40582] = 8'b1011101;
DRAM[40583] = 8'b1100110;
DRAM[40584] = 8'b1000110;
DRAM[40585] = 8'b101001;
DRAM[40586] = 8'b10000;
DRAM[40587] = 8'b1011;
DRAM[40588] = 8'b1100;
DRAM[40589] = 8'b111;
DRAM[40590] = 8'b11;
DRAM[40591] = 8'b11;
DRAM[40592] = 8'b11;
DRAM[40593] = 8'b10;
DRAM[40594] = 8'b0;
DRAM[40595] = 8'b1;
DRAM[40596] = 8'b11;
DRAM[40597] = 8'b100;
DRAM[40598] = 8'b11;
DRAM[40599] = 8'b10;
DRAM[40600] = 8'b0;
DRAM[40601] = 8'b1;
DRAM[40602] = 8'b0;
DRAM[40603] = 8'b101;
DRAM[40604] = 8'b1000;
DRAM[40605] = 8'b100;
DRAM[40606] = 8'b10010;
DRAM[40607] = 8'b110010;
DRAM[40608] = 8'b1100010;
DRAM[40609] = 8'b1110000;
DRAM[40610] = 8'b1010111;
DRAM[40611] = 8'b1011101;
DRAM[40612] = 8'b1111101;
DRAM[40613] = 8'b10010001;
DRAM[40614] = 8'b10101001;
DRAM[40615] = 8'b10101110;
DRAM[40616] = 8'b10111000;
DRAM[40617] = 8'b10111111;
DRAM[40618] = 8'b11001000;
DRAM[40619] = 8'b11001101;
DRAM[40620] = 8'b11010000;
DRAM[40621] = 8'b11010101;
DRAM[40622] = 8'b11011111;
DRAM[40623] = 8'b11100111;
DRAM[40624] = 8'b11101101;
DRAM[40625] = 8'b11101100;
DRAM[40626] = 8'b11100100;
DRAM[40627] = 8'b11011001;
DRAM[40628] = 8'b11010110;
DRAM[40629] = 8'b11011010;
DRAM[40630] = 8'b11011000;
DRAM[40631] = 8'b11010001;
DRAM[40632] = 8'b11001110;
DRAM[40633] = 8'b11010001;
DRAM[40634] = 8'b11001110;
DRAM[40635] = 8'b11000001;
DRAM[40636] = 8'b10110011;
DRAM[40637] = 8'b10101111;
DRAM[40638] = 8'b10111001;
DRAM[40639] = 8'b11000101;
DRAM[40640] = 8'b10111100;
DRAM[40641] = 8'b10111011;
DRAM[40642] = 8'b11000010;
DRAM[40643] = 8'b11001111;
DRAM[40644] = 8'b11010011;
DRAM[40645] = 8'b11001100;
DRAM[40646] = 8'b11001100;
DRAM[40647] = 8'b11010010;
DRAM[40648] = 8'b11010010;
DRAM[40649] = 8'b11000100;
DRAM[40650] = 8'b10110101;
DRAM[40651] = 8'b10110011;
DRAM[40652] = 8'b10111000;
DRAM[40653] = 8'b10110110;
DRAM[40654] = 8'b10101000;
DRAM[40655] = 8'b10011001;
DRAM[40656] = 8'b10011011;
DRAM[40657] = 8'b10011011;
DRAM[40658] = 8'b10011010;
DRAM[40659] = 8'b10011000;
DRAM[40660] = 8'b10010101;
DRAM[40661] = 8'b10010100;
DRAM[40662] = 8'b10010011;
DRAM[40663] = 8'b10010011;
DRAM[40664] = 8'b10010100;
DRAM[40665] = 8'b10010100;
DRAM[40666] = 8'b10010100;
DRAM[40667] = 8'b10010010;
DRAM[40668] = 8'b10001111;
DRAM[40669] = 8'b10001011;
DRAM[40670] = 8'b10001000;
DRAM[40671] = 8'b10000110;
DRAM[40672] = 8'b10001010;
DRAM[40673] = 8'b10001001;
DRAM[40674] = 8'b10000110;
DRAM[40675] = 8'b10000100;
DRAM[40676] = 8'b10000010;
DRAM[40677] = 8'b10000010;
DRAM[40678] = 8'b10000011;
DRAM[40679] = 8'b10000100;
DRAM[40680] = 8'b10000001;
DRAM[40681] = 8'b10000000;
DRAM[40682] = 8'b1111111;
DRAM[40683] = 8'b1111110;
DRAM[40684] = 8'b1111110;
DRAM[40685] = 8'b1111110;
DRAM[40686] = 8'b1111110;
DRAM[40687] = 8'b1111111;
DRAM[40688] = 8'b1111111;
DRAM[40689] = 8'b1111111;
DRAM[40690] = 8'b1111111;
DRAM[40691] = 8'b10000000;
DRAM[40692] = 8'b10000000;
DRAM[40693] = 8'b10000000;
DRAM[40694] = 8'b10000001;
DRAM[40695] = 8'b10000001;
DRAM[40696] = 8'b10000010;
DRAM[40697] = 8'b10000010;
DRAM[40698] = 8'b10000001;
DRAM[40699] = 8'b10000000;
DRAM[40700] = 8'b1111111;
DRAM[40701] = 8'b1111111;
DRAM[40702] = 8'b1111110;
DRAM[40703] = 8'b1111110;
DRAM[40704] = 8'b10011000;
DRAM[40705] = 8'b10011000;
DRAM[40706] = 8'b10011000;
DRAM[40707] = 8'b10011001;
DRAM[40708] = 8'b10011001;
DRAM[40709] = 8'b10011010;
DRAM[40710] = 8'b10011010;
DRAM[40711] = 8'b10011010;
DRAM[40712] = 8'b10011100;
DRAM[40713] = 8'b10011100;
DRAM[40714] = 8'b10011100;
DRAM[40715] = 8'b10011101;
DRAM[40716] = 8'b10011110;
DRAM[40717] = 8'b10011111;
DRAM[40718] = 8'b10100001;
DRAM[40719] = 8'b10100001;
DRAM[40720] = 8'b10011111;
DRAM[40721] = 8'b10011111;
DRAM[40722] = 8'b10100000;
DRAM[40723] = 8'b10100001;
DRAM[40724] = 8'b10100001;
DRAM[40725] = 8'b10100010;
DRAM[40726] = 8'b10100011;
DRAM[40727] = 8'b10100011;
DRAM[40728] = 8'b10100101;
DRAM[40729] = 8'b10100100;
DRAM[40730] = 8'b10100100;
DRAM[40731] = 8'b10100100;
DRAM[40732] = 8'b10100100;
DRAM[40733] = 8'b10100101;
DRAM[40734] = 8'b10100110;
DRAM[40735] = 8'b10100111;
DRAM[40736] = 8'b10100110;
DRAM[40737] = 8'b10100110;
DRAM[40738] = 8'b10100110;
DRAM[40739] = 8'b10100110;
DRAM[40740] = 8'b10100110;
DRAM[40741] = 8'b10100110;
DRAM[40742] = 8'b10100110;
DRAM[40743] = 8'b10100110;
DRAM[40744] = 8'b10100101;
DRAM[40745] = 8'b10100101;
DRAM[40746] = 8'b10101000;
DRAM[40747] = 8'b10101111;
DRAM[40748] = 8'b10111001;
DRAM[40749] = 8'b11001011;
DRAM[40750] = 8'b11100111;
DRAM[40751] = 8'b11111110;
DRAM[40752] = 8'b11111010;
DRAM[40753] = 8'b11111010;
DRAM[40754] = 8'b11111110;
DRAM[40755] = 8'b11111111;
DRAM[40756] = 8'b11111111;
DRAM[40757] = 8'b11111011;
DRAM[40758] = 8'b11111010;
DRAM[40759] = 8'b11111111;
DRAM[40760] = 8'b11111111;
DRAM[40761] = 8'b11111110;
DRAM[40762] = 8'b11111110;
DRAM[40763] = 8'b11111111;
DRAM[40764] = 8'b11111111;
DRAM[40765] = 8'b11111110;
DRAM[40766] = 8'b11111010;
DRAM[40767] = 8'b11110110;
DRAM[40768] = 8'b11110000;
DRAM[40769] = 8'b11100110;
DRAM[40770] = 8'b11011010;
DRAM[40771] = 8'b11010100;
DRAM[40772] = 8'b11010001;
DRAM[40773] = 8'b11001011;
DRAM[40774] = 8'b11000001;
DRAM[40775] = 8'b10111000;
DRAM[40776] = 8'b10110100;
DRAM[40777] = 8'b10101011;
DRAM[40778] = 8'b10100110;
DRAM[40779] = 8'b10100111;
DRAM[40780] = 8'b10100101;
DRAM[40781] = 8'b10011110;
DRAM[40782] = 8'b10011100;
DRAM[40783] = 8'b10011110;
DRAM[40784] = 8'b10011100;
DRAM[40785] = 8'b10011011;
DRAM[40786] = 8'b10100001;
DRAM[40787] = 8'b10101100;
DRAM[40788] = 8'b10110010;
DRAM[40789] = 8'b10101101;
DRAM[40790] = 8'b10100100;
DRAM[40791] = 8'b10011111;
DRAM[40792] = 8'b10100011;
DRAM[40793] = 8'b10100100;
DRAM[40794] = 8'b10101100;
DRAM[40795] = 8'b10110111;
DRAM[40796] = 8'b10111001;
DRAM[40797] = 8'b10110100;
DRAM[40798] = 8'b10110010;
DRAM[40799] = 8'b10110101;
DRAM[40800] = 8'b11000011;
DRAM[40801] = 8'b11000001;
DRAM[40802] = 8'b10111111;
DRAM[40803] = 8'b10111100;
DRAM[40804] = 8'b10111011;
DRAM[40805] = 8'b10111100;
DRAM[40806] = 8'b11000000;
DRAM[40807] = 8'b11000010;
DRAM[40808] = 8'b10110001;
DRAM[40809] = 8'b10111110;
DRAM[40810] = 8'b11001000;
DRAM[40811] = 8'b11001010;
DRAM[40812] = 8'b11001110;
DRAM[40813] = 8'b11011000;
DRAM[40814] = 8'b11011100;
DRAM[40815] = 8'b11011010;
DRAM[40816] = 8'b11010100;
DRAM[40817] = 8'b11010001;
DRAM[40818] = 8'b11010101;
DRAM[40819] = 8'b11011111;
DRAM[40820] = 8'b11011111;
DRAM[40821] = 8'b11010110;
DRAM[40822] = 8'b11010011;
DRAM[40823] = 8'b11010111;
DRAM[40824] = 8'b11001000;
DRAM[40825] = 8'b10111101;
DRAM[40826] = 8'b11000001;
DRAM[40827] = 8'b11000010;
DRAM[40828] = 8'b10111010;
DRAM[40829] = 8'b11000100;
DRAM[40830] = 8'b11001010;
DRAM[40831] = 8'b10111011;
DRAM[40832] = 8'b10110111;
DRAM[40833] = 8'b10101001;
DRAM[40834] = 8'b10010111;
DRAM[40835] = 8'b10000100;
DRAM[40836] = 8'b1010011;
DRAM[40837] = 8'b111101;
DRAM[40838] = 8'b1011001;
DRAM[40839] = 8'b1011111;
DRAM[40840] = 8'b1000110;
DRAM[40841] = 8'b100010;
DRAM[40842] = 8'b1;
DRAM[40843] = 8'b0;
DRAM[40844] = 8'b100;
DRAM[40845] = 8'b100;
DRAM[40846] = 8'b1;
DRAM[40847] = 8'b1;
DRAM[40848] = 8'b0;
DRAM[40849] = 8'b0;
DRAM[40850] = 8'b0;
DRAM[40851] = 8'b0;
DRAM[40852] = 8'b1;
DRAM[40853] = 8'b10;
DRAM[40854] = 8'b10;
DRAM[40855] = 8'b0;
DRAM[40856] = 8'b0;
DRAM[40857] = 8'b0;
DRAM[40858] = 8'b0;
DRAM[40859] = 8'b111;
DRAM[40860] = 8'b1101;
DRAM[40861] = 8'b111;
DRAM[40862] = 8'b10011;
DRAM[40863] = 8'b110000;
DRAM[40864] = 8'b1010100;
DRAM[40865] = 8'b1100100;
DRAM[40866] = 8'b1010000;
DRAM[40867] = 8'b1100101;
DRAM[40868] = 8'b10001111;
DRAM[40869] = 8'b10011100;
DRAM[40870] = 8'b10101100;
DRAM[40871] = 8'b10101100;
DRAM[40872] = 8'b10110101;
DRAM[40873] = 8'b10111001;
DRAM[40874] = 8'b11000010;
DRAM[40875] = 8'b11001110;
DRAM[40876] = 8'b11011010;
DRAM[40877] = 8'b11100100;
DRAM[40878] = 8'b11101011;
DRAM[40879] = 8'b11101110;
DRAM[40880] = 8'b11101011;
DRAM[40881] = 8'b11101111;
DRAM[40882] = 8'b11100110;
DRAM[40883] = 8'b11010011;
DRAM[40884] = 8'b11001101;
DRAM[40885] = 8'b11010100;
DRAM[40886] = 8'b11010101;
DRAM[40887] = 8'b11001100;
DRAM[40888] = 8'b11000111;
DRAM[40889] = 8'b11010000;
DRAM[40890] = 8'b11010100;
DRAM[40891] = 8'b11001010;
DRAM[40892] = 8'b10111010;
DRAM[40893] = 8'b10110011;
DRAM[40894] = 8'b10111011;
DRAM[40895] = 8'b11000111;
DRAM[40896] = 8'b11001101;
DRAM[40897] = 8'b11001101;
DRAM[40898] = 8'b11010011;
DRAM[40899] = 8'b11011010;
DRAM[40900] = 8'b11010011;
DRAM[40901] = 8'b11000011;
DRAM[40902] = 8'b11000000;
DRAM[40903] = 8'b11001000;
DRAM[40904] = 8'b11010100;
DRAM[40905] = 8'b11001111;
DRAM[40906] = 8'b11000110;
DRAM[40907] = 8'b10111001;
DRAM[40908] = 8'b10101101;
DRAM[40909] = 8'b10100110;
DRAM[40910] = 8'b10100101;
DRAM[40911] = 8'b10100111;
DRAM[40912] = 8'b10011111;
DRAM[40913] = 8'b10011111;
DRAM[40914] = 8'b10011101;
DRAM[40915] = 8'b10011010;
DRAM[40916] = 8'b10010101;
DRAM[40917] = 8'b10010010;
DRAM[40918] = 8'b10010000;
DRAM[40919] = 8'b10010000;
DRAM[40920] = 8'b10010000;
DRAM[40921] = 8'b10010000;
DRAM[40922] = 8'b10001111;
DRAM[40923] = 8'b10001110;
DRAM[40924] = 8'b10001101;
DRAM[40925] = 8'b10001100;
DRAM[40926] = 8'b10001100;
DRAM[40927] = 8'b10001100;
DRAM[40928] = 8'b10001010;
DRAM[40929] = 8'b10001001;
DRAM[40930] = 8'b10000110;
DRAM[40931] = 8'b10000011;
DRAM[40932] = 8'b10000010;
DRAM[40933] = 8'b10000010;
DRAM[40934] = 8'b10000011;
DRAM[40935] = 8'b10000100;
DRAM[40936] = 8'b10000001;
DRAM[40937] = 8'b10000000;
DRAM[40938] = 8'b1111111;
DRAM[40939] = 8'b1111110;
DRAM[40940] = 8'b1111110;
DRAM[40941] = 8'b1111110;
DRAM[40942] = 8'b1111110;
DRAM[40943] = 8'b1111111;
DRAM[40944] = 8'b1111111;
DRAM[40945] = 8'b1111111;
DRAM[40946] = 8'b1111111;
DRAM[40947] = 8'b10000000;
DRAM[40948] = 8'b10000000;
DRAM[40949] = 8'b10000001;
DRAM[40950] = 8'b10000001;
DRAM[40951] = 8'b10000001;
DRAM[40952] = 8'b10000010;
DRAM[40953] = 8'b10000010;
DRAM[40954] = 8'b10000001;
DRAM[40955] = 8'b10000000;
DRAM[40956] = 8'b10000000;
DRAM[40957] = 8'b1111111;
DRAM[40958] = 8'b1111110;
DRAM[40959] = 8'b1111110;
DRAM[40960] = 8'b10010110;
DRAM[40961] = 8'b10010110;
DRAM[40962] = 8'b10010111;
DRAM[40963] = 8'b10011000;
DRAM[40964] = 8'b10011000;
DRAM[40965] = 8'b10011001;
DRAM[40966] = 8'b10011010;
DRAM[40967] = 8'b10011010;
DRAM[40968] = 8'b10011001;
DRAM[40969] = 8'b10011011;
DRAM[40970] = 8'b10011101;
DRAM[40971] = 8'b10011111;
DRAM[40972] = 8'b10100001;
DRAM[40973] = 8'b10100010;
DRAM[40974] = 8'b10100011;
DRAM[40975] = 8'b10100011;
DRAM[40976] = 8'b10011111;
DRAM[40977] = 8'b10011111;
DRAM[40978] = 8'b10100000;
DRAM[40979] = 8'b10100001;
DRAM[40980] = 8'b10100011;
DRAM[40981] = 8'b10100100;
DRAM[40982] = 8'b10100101;
DRAM[40983] = 8'b10100110;
DRAM[40984] = 8'b10100101;
DRAM[40985] = 8'b10100101;
DRAM[40986] = 8'b10100101;
DRAM[40987] = 8'b10100101;
DRAM[40988] = 8'b10100101;
DRAM[40989] = 8'b10100101;
DRAM[40990] = 8'b10100101;
DRAM[40991] = 8'b10100101;
DRAM[40992] = 8'b10100010;
DRAM[40993] = 8'b10100100;
DRAM[40994] = 8'b10100110;
DRAM[40995] = 8'b10100110;
DRAM[40996] = 8'b10100110;
DRAM[40997] = 8'b10100101;
DRAM[40998] = 8'b10100101;
DRAM[40999] = 8'b10100110;
DRAM[41000] = 8'b10101001;
DRAM[41001] = 8'b10100011;
DRAM[41002] = 8'b10100100;
DRAM[41003] = 8'b10110100;
DRAM[41004] = 8'b11001111;
DRAM[41005] = 8'b11101001;
DRAM[41006] = 8'b11111100;
DRAM[41007] = 8'b11111111;
DRAM[41008] = 8'b11111110;
DRAM[41009] = 8'b11111110;
DRAM[41010] = 8'b11111110;
DRAM[41011] = 8'b11111110;
DRAM[41012] = 8'b11111110;
DRAM[41013] = 8'b11111110;
DRAM[41014] = 8'b11111110;
DRAM[41015] = 8'b11111110;
DRAM[41016] = 8'b11111110;
DRAM[41017] = 8'b11111101;
DRAM[41018] = 8'b11111101;
DRAM[41019] = 8'b11111110;
DRAM[41020] = 8'b11111111;
DRAM[41021] = 8'b11111110;
DRAM[41022] = 8'b11111100;
DRAM[41023] = 8'b11111001;
DRAM[41024] = 8'b11110000;
DRAM[41025] = 8'b11101001;
DRAM[41026] = 8'b11100000;
DRAM[41027] = 8'b11011001;
DRAM[41028] = 8'b11010100;
DRAM[41029] = 8'b11001101;
DRAM[41030] = 8'b11000101;
DRAM[41031] = 8'b11000000;
DRAM[41032] = 8'b10111100;
DRAM[41033] = 8'b10110101;
DRAM[41034] = 8'b10101010;
DRAM[41035] = 8'b10100010;
DRAM[41036] = 8'b10100011;
DRAM[41037] = 8'b10100111;
DRAM[41038] = 8'b10100101;
DRAM[41039] = 8'b10011111;
DRAM[41040] = 8'b10011000;
DRAM[41041] = 8'b10011001;
DRAM[41042] = 8'b10011100;
DRAM[41043] = 8'b10100001;
DRAM[41044] = 8'b10100100;
DRAM[41045] = 8'b10100100;
DRAM[41046] = 8'b10100000;
DRAM[41047] = 8'b10011101;
DRAM[41048] = 8'b10011001;
DRAM[41049] = 8'b10100101;
DRAM[41050] = 8'b10110010;
DRAM[41051] = 8'b10110100;
DRAM[41052] = 8'b10101101;
DRAM[41053] = 8'b10100111;
DRAM[41054] = 8'b10100111;
DRAM[41055] = 8'b10101011;
DRAM[41056] = 8'b10110101;
DRAM[41057] = 8'b10110111;
DRAM[41058] = 8'b10111001;
DRAM[41059] = 8'b10111010;
DRAM[41060] = 8'b10111001;
DRAM[41061] = 8'b10111000;
DRAM[41062] = 8'b10111000;
DRAM[41063] = 8'b10111001;
DRAM[41064] = 8'b10111010;
DRAM[41065] = 8'b11000011;
DRAM[41066] = 8'b11001101;
DRAM[41067] = 8'b11010101;
DRAM[41068] = 8'b11010111;
DRAM[41069] = 8'b11010111;
DRAM[41070] = 8'b11011001;
DRAM[41071] = 8'b11011010;
DRAM[41072] = 8'b11001100;
DRAM[41073] = 8'b11010001;
DRAM[41074] = 8'b11011100;
DRAM[41075] = 8'b11011101;
DRAM[41076] = 8'b11010011;
DRAM[41077] = 8'b11010001;
DRAM[41078] = 8'b11010000;
DRAM[41079] = 8'b11000110;
DRAM[41080] = 8'b10111000;
DRAM[41081] = 8'b10110010;
DRAM[41082] = 8'b10101100;
DRAM[41083] = 8'b10101110;
DRAM[41084] = 8'b10110101;
DRAM[41085] = 8'b10111110;
DRAM[41086] = 8'b11000011;
DRAM[41087] = 8'b11000101;
DRAM[41088] = 8'b11000010;
DRAM[41089] = 8'b10101010;
DRAM[41090] = 8'b10010000;
DRAM[41091] = 8'b1111001;
DRAM[41092] = 8'b1011011;
DRAM[41093] = 8'b1000010;
DRAM[41094] = 8'b1001001;
DRAM[41095] = 8'b1100000;
DRAM[41096] = 8'b1000001;
DRAM[41097] = 8'b11010;
DRAM[41098] = 8'b100;
DRAM[41099] = 8'b100;
DRAM[41100] = 8'b11;
DRAM[41101] = 8'b11;
DRAM[41102] = 8'b101;
DRAM[41103] = 8'b11;
DRAM[41104] = 8'b0;
DRAM[41105] = 8'b0;
DRAM[41106] = 8'b0;
DRAM[41107] = 8'b0;
DRAM[41108] = 8'b0;
DRAM[41109] = 8'b0;
DRAM[41110] = 8'b0;
DRAM[41111] = 8'b0;
DRAM[41112] = 8'b0;
DRAM[41113] = 8'b0;
DRAM[41114] = 8'b1;
DRAM[41115] = 8'b11;
DRAM[41116] = 8'b1010;
DRAM[41117] = 8'b11010;
DRAM[41118] = 8'b101111;
DRAM[41119] = 8'b111111;
DRAM[41120] = 8'b1010111;
DRAM[41121] = 8'b1001000;
DRAM[41122] = 8'b1001100;
DRAM[41123] = 8'b1100110;
DRAM[41124] = 8'b10000111;
DRAM[41125] = 8'b10100100;
DRAM[41126] = 8'b10101110;
DRAM[41127] = 8'b10100101;
DRAM[41128] = 8'b10011011;
DRAM[41129] = 8'b10100110;
DRAM[41130] = 8'b10111011;
DRAM[41131] = 8'b11010001;
DRAM[41132] = 8'b11011110;
DRAM[41133] = 8'b11100100;
DRAM[41134] = 8'b11101010;
DRAM[41135] = 8'b11110000;
DRAM[41136] = 8'b11101111;
DRAM[41137] = 8'b11110100;
DRAM[41138] = 8'b11110100;
DRAM[41139] = 8'b11101001;
DRAM[41140] = 8'b11011010;
DRAM[41141] = 8'b11010000;
DRAM[41142] = 8'b11001111;
DRAM[41143] = 8'b11010000;
DRAM[41144] = 8'b11010101;
DRAM[41145] = 8'b11010011;
DRAM[41146] = 8'b11010110;
DRAM[41147] = 8'b10111111;
DRAM[41148] = 8'b10110011;
DRAM[41149] = 8'b10111000;
DRAM[41150] = 8'b10110000;
DRAM[41151] = 8'b10110011;
DRAM[41152] = 8'b10110111;
DRAM[41153] = 8'b11000110;
DRAM[41154] = 8'b11010100;
DRAM[41155] = 8'b11011110;
DRAM[41156] = 8'b11101001;
DRAM[41157] = 8'b11101011;
DRAM[41158] = 8'b11011000;
DRAM[41159] = 8'b11000000;
DRAM[41160] = 8'b10110111;
DRAM[41161] = 8'b10111001;
DRAM[41162] = 8'b10111001;
DRAM[41163] = 8'b10110101;
DRAM[41164] = 8'b10101110;
DRAM[41165] = 8'b10100101;
DRAM[41166] = 8'b10011111;
DRAM[41167] = 8'b10011100;
DRAM[41168] = 8'b10100011;
DRAM[41169] = 8'b10100000;
DRAM[41170] = 8'b10011101;
DRAM[41171] = 8'b10011011;
DRAM[41172] = 8'b10011010;
DRAM[41173] = 8'b10011001;
DRAM[41174] = 8'b10010111;
DRAM[41175] = 8'b10010101;
DRAM[41176] = 8'b10010101;
DRAM[41177] = 8'b10010011;
DRAM[41178] = 8'b10010001;
DRAM[41179] = 8'b10001111;
DRAM[41180] = 8'b10001101;
DRAM[41181] = 8'b10001100;
DRAM[41182] = 8'b10001011;
DRAM[41183] = 8'b10001011;
DRAM[41184] = 8'b10001100;
DRAM[41185] = 8'b10001000;
DRAM[41186] = 8'b10000100;
DRAM[41187] = 8'b10000010;
DRAM[41188] = 8'b10000011;
DRAM[41189] = 8'b10000100;
DRAM[41190] = 8'b10000100;
DRAM[41191] = 8'b10000011;
DRAM[41192] = 8'b10000001;
DRAM[41193] = 8'b10000000;
DRAM[41194] = 8'b1111111;
DRAM[41195] = 8'b1111110;
DRAM[41196] = 8'b1111101;
DRAM[41197] = 8'b1111100;
DRAM[41198] = 8'b1111100;
DRAM[41199] = 8'b1111100;
DRAM[41200] = 8'b1111010;
DRAM[41201] = 8'b1111100;
DRAM[41202] = 8'b1111111;
DRAM[41203] = 8'b10000010;
DRAM[41204] = 8'b10000011;
DRAM[41205] = 8'b10000011;
DRAM[41206] = 8'b10000010;
DRAM[41207] = 8'b10000001;
DRAM[41208] = 8'b10000101;
DRAM[41209] = 8'b10000010;
DRAM[41210] = 8'b1111111;
DRAM[41211] = 8'b1111111;
DRAM[41212] = 8'b10000000;
DRAM[41213] = 8'b10000001;
DRAM[41214] = 8'b10000001;
DRAM[41215] = 8'b10000000;
DRAM[41216] = 8'b10010110;
DRAM[41217] = 8'b10010110;
DRAM[41218] = 8'b10010111;
DRAM[41219] = 8'b10011000;
DRAM[41220] = 8'b10011000;
DRAM[41221] = 8'b10011001;
DRAM[41222] = 8'b10011010;
DRAM[41223] = 8'b10011010;
DRAM[41224] = 8'b10011010;
DRAM[41225] = 8'b10011011;
DRAM[41226] = 8'b10011101;
DRAM[41227] = 8'b10011111;
DRAM[41228] = 8'b10100000;
DRAM[41229] = 8'b10100001;
DRAM[41230] = 8'b10100010;
DRAM[41231] = 8'b10100010;
DRAM[41232] = 8'b10011101;
DRAM[41233] = 8'b10011110;
DRAM[41234] = 8'b10011111;
DRAM[41235] = 8'b10100000;
DRAM[41236] = 8'b10100001;
DRAM[41237] = 8'b10100011;
DRAM[41238] = 8'b10100100;
DRAM[41239] = 8'b10100100;
DRAM[41240] = 8'b10100101;
DRAM[41241] = 8'b10100101;
DRAM[41242] = 8'b10100101;
DRAM[41243] = 8'b10100101;
DRAM[41244] = 8'b10100101;
DRAM[41245] = 8'b10100101;
DRAM[41246] = 8'b10100101;
DRAM[41247] = 8'b10100101;
DRAM[41248] = 8'b10101010;
DRAM[41249] = 8'b10101001;
DRAM[41250] = 8'b10100111;
DRAM[41251] = 8'b10100110;
DRAM[41252] = 8'b10100101;
DRAM[41253] = 8'b10100101;
DRAM[41254] = 8'b10100101;
DRAM[41255] = 8'b10100101;
DRAM[41256] = 8'b10101010;
DRAM[41257] = 8'b10101010;
DRAM[41258] = 8'b10110001;
DRAM[41259] = 8'b11000101;
DRAM[41260] = 8'b11011111;
DRAM[41261] = 8'b11110011;
DRAM[41262] = 8'b11111101;
DRAM[41263] = 8'b11111111;
DRAM[41264] = 8'b11111110;
DRAM[41265] = 8'b11111110;
DRAM[41266] = 8'b11111110;
DRAM[41267] = 8'b11111110;
DRAM[41268] = 8'b11111110;
DRAM[41269] = 8'b11111110;
DRAM[41270] = 8'b11111110;
DRAM[41271] = 8'b11111110;
DRAM[41272] = 8'b11111110;
DRAM[41273] = 8'b11111101;
DRAM[41274] = 8'b11111101;
DRAM[41275] = 8'b11111110;
DRAM[41276] = 8'b11111111;
DRAM[41277] = 8'b11111110;
DRAM[41278] = 8'b11111011;
DRAM[41279] = 8'b11111000;
DRAM[41280] = 8'b11110001;
DRAM[41281] = 8'b11101010;
DRAM[41282] = 8'b11100000;
DRAM[41283] = 8'b11011001;
DRAM[41284] = 8'b11010100;
DRAM[41285] = 8'b11001110;
DRAM[41286] = 8'b11001000;
DRAM[41287] = 8'b11000011;
DRAM[41288] = 8'b10111111;
DRAM[41289] = 8'b10111110;
DRAM[41290] = 8'b10111001;
DRAM[41291] = 8'b10110000;
DRAM[41292] = 8'b10101001;
DRAM[41293] = 8'b10100110;
DRAM[41294] = 8'b10100000;
DRAM[41295] = 8'b10011010;
DRAM[41296] = 8'b10010100;
DRAM[41297] = 8'b10010101;
DRAM[41298] = 8'b10011000;
DRAM[41299] = 8'b10011101;
DRAM[41300] = 8'b10100010;
DRAM[41301] = 8'b10100100;
DRAM[41302] = 8'b10100011;
DRAM[41303] = 8'b10100001;
DRAM[41304] = 8'b10101010;
DRAM[41305] = 8'b10101100;
DRAM[41306] = 8'b10101101;
DRAM[41307] = 8'b10101101;
DRAM[41308] = 8'b10101011;
DRAM[41309] = 8'b10101011;
DRAM[41310] = 8'b10101110;
DRAM[41311] = 8'b10110000;
DRAM[41312] = 8'b10101011;
DRAM[41313] = 8'b10110001;
DRAM[41314] = 8'b10111000;
DRAM[41315] = 8'b10111101;
DRAM[41316] = 8'b10111110;
DRAM[41317] = 8'b10111100;
DRAM[41318] = 8'b10111010;
DRAM[41319] = 8'b10111001;
DRAM[41320] = 8'b11000101;
DRAM[41321] = 8'b11001001;
DRAM[41322] = 8'b11001111;
DRAM[41323] = 8'b11010011;
DRAM[41324] = 8'b11010011;
DRAM[41325] = 8'b11010010;
DRAM[41326] = 8'b11010001;
DRAM[41327] = 8'b11010000;
DRAM[41328] = 8'b11001011;
DRAM[41329] = 8'b11001001;
DRAM[41330] = 8'b11010000;
DRAM[41331] = 8'b11010100;
DRAM[41332] = 8'b11010001;
DRAM[41333] = 8'b11010000;
DRAM[41334] = 8'b11000111;
DRAM[41335] = 8'b10110100;
DRAM[41336] = 8'b10101010;
DRAM[41337] = 8'b10101001;
DRAM[41338] = 8'b10100101;
DRAM[41339] = 8'b10100001;
DRAM[41340] = 8'b10100101;
DRAM[41341] = 8'b10110010;
DRAM[41342] = 8'b10111100;
DRAM[41343] = 8'b11000000;
DRAM[41344] = 8'b10110110;
DRAM[41345] = 8'b10101010;
DRAM[41346] = 8'b10011001;
DRAM[41347] = 8'b1111101;
DRAM[41348] = 8'b1010011;
DRAM[41349] = 8'b110011;
DRAM[41350] = 8'b111011;
DRAM[41351] = 8'b1010101;
DRAM[41352] = 8'b110101;
DRAM[41353] = 8'b11101;
DRAM[41354] = 8'b1111;
DRAM[41355] = 8'b1011;
DRAM[41356] = 8'b1;
DRAM[41357] = 8'b0;
DRAM[41358] = 8'b1;
DRAM[41359] = 8'b0;
DRAM[41360] = 8'b0;
DRAM[41361] = 8'b0;
DRAM[41362] = 8'b0;
DRAM[41363] = 8'b0;
DRAM[41364] = 8'b0;
DRAM[41365] = 8'b0;
DRAM[41366] = 8'b0;
DRAM[41367] = 8'b0;
DRAM[41368] = 8'b11;
DRAM[41369] = 8'b100;
DRAM[41370] = 8'b100;
DRAM[41371] = 8'b101;
DRAM[41372] = 8'b1010;
DRAM[41373] = 8'b10110;
DRAM[41374] = 8'b100111;
DRAM[41375] = 8'b110100;
DRAM[41376] = 8'b111010;
DRAM[41377] = 8'b111100;
DRAM[41378] = 8'b1001100;
DRAM[41379] = 8'b1110000;
DRAM[41380] = 8'b10010101;
DRAM[41381] = 8'b10100111;
DRAM[41382] = 8'b10101000;
DRAM[41383] = 8'b10101000;
DRAM[41384] = 8'b10001111;
DRAM[41385] = 8'b10011001;
DRAM[41386] = 8'b10101011;
DRAM[41387] = 8'b11000000;
DRAM[41388] = 8'b11001111;
DRAM[41389] = 8'b11010111;
DRAM[41390] = 8'b11100001;
DRAM[41391] = 8'b11101011;
DRAM[41392] = 8'b11101000;
DRAM[41393] = 8'b11101100;
DRAM[41394] = 8'b11101011;
DRAM[41395] = 8'b11100100;
DRAM[41396] = 8'b11011101;
DRAM[41397] = 8'b11011010;
DRAM[41398] = 8'b11011010;
DRAM[41399] = 8'b11011001;
DRAM[41400] = 8'b11010000;
DRAM[41401] = 8'b11011001;
DRAM[41402] = 8'b11100110;
DRAM[41403] = 8'b11001111;
DRAM[41404] = 8'b10111100;
DRAM[41405] = 8'b10111111;
DRAM[41406] = 8'b10111101;
DRAM[41407] = 8'b11001000;
DRAM[41408] = 8'b11000101;
DRAM[41409] = 8'b11010001;
DRAM[41410] = 8'b11010010;
DRAM[41411] = 8'b11000100;
DRAM[41412] = 8'b10111011;
DRAM[41413] = 8'b11000111;
DRAM[41414] = 8'b11011010;
DRAM[41415] = 8'b11100100;
DRAM[41416] = 8'b11101010;
DRAM[41417] = 8'b11011111;
DRAM[41418] = 8'b11001100;
DRAM[41419] = 8'b10110110;
DRAM[41420] = 8'b10100100;
DRAM[41421] = 8'b10011110;
DRAM[41422] = 8'b10100000;
DRAM[41423] = 8'b10100101;
DRAM[41424] = 8'b10011110;
DRAM[41425] = 8'b10011111;
DRAM[41426] = 8'b10100001;
DRAM[41427] = 8'b10100010;
DRAM[41428] = 8'b10100001;
DRAM[41429] = 8'b10011010;
DRAM[41430] = 8'b10010001;
DRAM[41431] = 8'b10001011;
DRAM[41432] = 8'b10010000;
DRAM[41433] = 8'b10010000;
DRAM[41434] = 8'b10001111;
DRAM[41435] = 8'b10001111;
DRAM[41436] = 8'b10001110;
DRAM[41437] = 8'b10001110;
DRAM[41438] = 8'b10001111;
DRAM[41439] = 8'b10001111;
DRAM[41440] = 8'b10001100;
DRAM[41441] = 8'b10001001;
DRAM[41442] = 8'b10000101;
DRAM[41443] = 8'b10000100;
DRAM[41444] = 8'b10000100;
DRAM[41445] = 8'b10000101;
DRAM[41446] = 8'b10000101;
DRAM[41447] = 8'b10000100;
DRAM[41448] = 8'b10000001;
DRAM[41449] = 8'b10000000;
DRAM[41450] = 8'b1111111;
DRAM[41451] = 8'b1111110;
DRAM[41452] = 8'b1111101;
DRAM[41453] = 8'b1111100;
DRAM[41454] = 8'b1111100;
DRAM[41455] = 8'b1111100;
DRAM[41456] = 8'b1111011;
DRAM[41457] = 8'b1111101;
DRAM[41458] = 8'b1111111;
DRAM[41459] = 8'b10000010;
DRAM[41460] = 8'b10000011;
DRAM[41461] = 8'b10000011;
DRAM[41462] = 8'b10000010;
DRAM[41463] = 8'b10000001;
DRAM[41464] = 8'b10000101;
DRAM[41465] = 8'b10000011;
DRAM[41466] = 8'b10000000;
DRAM[41467] = 8'b1111111;
DRAM[41468] = 8'b10000000;
DRAM[41469] = 8'b10000001;
DRAM[41470] = 8'b10000001;
DRAM[41471] = 8'b10000000;
DRAM[41472] = 8'b10010110;
DRAM[41473] = 8'b10010110;
DRAM[41474] = 8'b10010111;
DRAM[41475] = 8'b10011000;
DRAM[41476] = 8'b10011000;
DRAM[41477] = 8'b10011001;
DRAM[41478] = 8'b10011010;
DRAM[41479] = 8'b10011010;
DRAM[41480] = 8'b10011011;
DRAM[41481] = 8'b10011100;
DRAM[41482] = 8'b10011110;
DRAM[41483] = 8'b10011111;
DRAM[41484] = 8'b10100000;
DRAM[41485] = 8'b10100000;
DRAM[41486] = 8'b10100000;
DRAM[41487] = 8'b10100000;
DRAM[41488] = 8'b10011101;
DRAM[41489] = 8'b10011101;
DRAM[41490] = 8'b10011110;
DRAM[41491] = 8'b10011111;
DRAM[41492] = 8'b10100000;
DRAM[41493] = 8'b10100001;
DRAM[41494] = 8'b10100010;
DRAM[41495] = 8'b10100011;
DRAM[41496] = 8'b10100100;
DRAM[41497] = 8'b10100100;
DRAM[41498] = 8'b10100100;
DRAM[41499] = 8'b10100101;
DRAM[41500] = 8'b10100101;
DRAM[41501] = 8'b10100101;
DRAM[41502] = 8'b10100101;
DRAM[41503] = 8'b10100101;
DRAM[41504] = 8'b10101010;
DRAM[41505] = 8'b10100111;
DRAM[41506] = 8'b10100011;
DRAM[41507] = 8'b10100001;
DRAM[41508] = 8'b10100010;
DRAM[41509] = 8'b10100100;
DRAM[41510] = 8'b10100101;
DRAM[41511] = 8'b10100110;
DRAM[41512] = 8'b10101100;
DRAM[41513] = 8'b10110111;
DRAM[41514] = 8'b11001001;
DRAM[41515] = 8'b11011111;
DRAM[41516] = 8'b11110010;
DRAM[41517] = 8'b11111101;
DRAM[41518] = 8'b11111101;
DRAM[41519] = 8'b11111010;
DRAM[41520] = 8'b11111110;
DRAM[41521] = 8'b11111110;
DRAM[41522] = 8'b11111110;
DRAM[41523] = 8'b11111110;
DRAM[41524] = 8'b11111110;
DRAM[41525] = 8'b11111110;
DRAM[41526] = 8'b11111110;
DRAM[41527] = 8'b11111110;
DRAM[41528] = 8'b11111110;
DRAM[41529] = 8'b11111101;
DRAM[41530] = 8'b11111101;
DRAM[41531] = 8'b11111110;
DRAM[41532] = 8'b11111110;
DRAM[41533] = 8'b11111101;
DRAM[41534] = 8'b11111010;
DRAM[41535] = 8'b11110111;
DRAM[41536] = 8'b11110001;
DRAM[41537] = 8'b11101001;
DRAM[41538] = 8'b11011111;
DRAM[41539] = 8'b11010111;
DRAM[41540] = 8'b11010011;
DRAM[41541] = 8'b11001111;
DRAM[41542] = 8'b11001010;
DRAM[41543] = 8'b11000110;
DRAM[41544] = 8'b10111101;
DRAM[41545] = 8'b10111111;
DRAM[41546] = 8'b10111011;
DRAM[41547] = 8'b10101111;
DRAM[41548] = 8'b10100101;
DRAM[41549] = 8'b10100000;
DRAM[41550] = 8'b10011100;
DRAM[41551] = 8'b10011000;
DRAM[41552] = 8'b10010111;
DRAM[41553] = 8'b10010111;
DRAM[41554] = 8'b10010111;
DRAM[41555] = 8'b10011011;
DRAM[41556] = 8'b10011111;
DRAM[41557] = 8'b10100010;
DRAM[41558] = 8'b10100010;
DRAM[41559] = 8'b10100001;
DRAM[41560] = 8'b10100001;
DRAM[41561] = 8'b10100011;
DRAM[41562] = 8'b10101001;
DRAM[41563] = 8'b10110001;
DRAM[41564] = 8'b10110111;
DRAM[41565] = 8'b10110101;
DRAM[41566] = 8'b10101110;
DRAM[41567] = 8'b10100110;
DRAM[41568] = 8'b10100011;
DRAM[41569] = 8'b10101000;
DRAM[41570] = 8'b10110000;
DRAM[41571] = 8'b10110110;
DRAM[41572] = 8'b10111001;
DRAM[41573] = 8'b10111010;
DRAM[41574] = 8'b10111011;
DRAM[41575] = 8'b10111100;
DRAM[41576] = 8'b11000101;
DRAM[41577] = 8'b11000111;
DRAM[41578] = 8'b11001010;
DRAM[41579] = 8'b11001110;
DRAM[41580] = 8'b11010010;
DRAM[41581] = 8'b11010011;
DRAM[41582] = 8'b11010010;
DRAM[41583] = 8'b11010000;
DRAM[41584] = 8'b11001110;
DRAM[41585] = 8'b11001000;
DRAM[41586] = 8'b11001100;
DRAM[41587] = 8'b11010100;
DRAM[41588] = 8'b11010110;
DRAM[41589] = 8'b11010111;
DRAM[41590] = 8'b11001011;
DRAM[41591] = 8'b10110011;
DRAM[41592] = 8'b10100110;
DRAM[41593] = 8'b10101101;
DRAM[41594] = 8'b10101001;
DRAM[41595] = 8'b10011101;
DRAM[41596] = 8'b10011110;
DRAM[41597] = 8'b10101101;
DRAM[41598] = 8'b10111000;
DRAM[41599] = 8'b10111000;
DRAM[41600] = 8'b10101110;
DRAM[41601] = 8'b10100111;
DRAM[41602] = 8'b10011011;
DRAM[41603] = 8'b10000010;
DRAM[41604] = 8'b1011001;
DRAM[41605] = 8'b110100;
DRAM[41606] = 8'b101111;
DRAM[41607] = 8'b111101;
DRAM[41608] = 8'b101100;
DRAM[41609] = 8'b100011;
DRAM[41610] = 8'b100000;
DRAM[41611] = 8'b10110;
DRAM[41612] = 8'b100;
DRAM[41613] = 8'b0;
DRAM[41614] = 8'b11;
DRAM[41615] = 8'b0;
DRAM[41616] = 8'b0;
DRAM[41617] = 8'b0;
DRAM[41618] = 8'b0;
DRAM[41619] = 8'b0;
DRAM[41620] = 8'b0;
DRAM[41621] = 8'b0;
DRAM[41622] = 8'b0;
DRAM[41623] = 8'b0;
DRAM[41624] = 8'b1;
DRAM[41625] = 8'b1;
DRAM[41626] = 8'b1;
DRAM[41627] = 8'b1;
DRAM[41628] = 8'b11;
DRAM[41629] = 8'b1010;
DRAM[41630] = 8'b10110;
DRAM[41631] = 8'b11111;
DRAM[41632] = 8'b100010;
DRAM[41633] = 8'b110110;
DRAM[41634] = 8'b1001100;
DRAM[41635] = 8'b1110011;
DRAM[41636] = 8'b10011001;
DRAM[41637] = 8'b10011011;
DRAM[41638] = 8'b10010110;
DRAM[41639] = 8'b10100111;
DRAM[41640] = 8'b10011101;
DRAM[41641] = 8'b10100010;
DRAM[41642] = 8'b10101110;
DRAM[41643] = 8'b10111100;
DRAM[41644] = 8'b11000111;
DRAM[41645] = 8'b11010000;
DRAM[41646] = 8'b11011100;
DRAM[41647] = 8'b11101000;
DRAM[41648] = 8'b11100100;
DRAM[41649] = 8'b11100111;
DRAM[41650] = 8'b11100110;
DRAM[41651] = 8'b11100000;
DRAM[41652] = 8'b11011110;
DRAM[41653] = 8'b11100000;
DRAM[41654] = 8'b11100000;
DRAM[41655] = 8'b11011101;
DRAM[41656] = 8'b11001011;
DRAM[41657] = 8'b11010010;
DRAM[41658] = 8'b11011110;
DRAM[41659] = 8'b11001000;
DRAM[41660] = 8'b10110111;
DRAM[41661] = 8'b10111010;
DRAM[41662] = 8'b10110100;
DRAM[41663] = 8'b10111100;
DRAM[41664] = 8'b10110111;
DRAM[41665] = 8'b11000110;
DRAM[41666] = 8'b11010010;
DRAM[41667] = 8'b11010010;
DRAM[41668] = 8'b11001111;
DRAM[41669] = 8'b11001101;
DRAM[41670] = 8'b11000111;
DRAM[41671] = 8'b10111111;
DRAM[41672] = 8'b10111100;
DRAM[41673] = 8'b11000110;
DRAM[41674] = 8'b11010010;
DRAM[41675] = 8'b11010110;
DRAM[41676] = 8'b11001101;
DRAM[41677] = 8'b10111011;
DRAM[41678] = 8'b10100110;
DRAM[41679] = 8'b10011010;
DRAM[41680] = 8'b10011011;
DRAM[41681] = 8'b10011000;
DRAM[41682] = 8'b10010101;
DRAM[41683] = 8'b10010101;
DRAM[41684] = 8'b10011000;
DRAM[41685] = 8'b10011011;
DRAM[41686] = 8'b10011101;
DRAM[41687] = 8'b10011110;
DRAM[41688] = 8'b10010101;
DRAM[41689] = 8'b10010100;
DRAM[41690] = 8'b10010010;
DRAM[41691] = 8'b10010000;
DRAM[41692] = 8'b10001110;
DRAM[41693] = 8'b10001100;
DRAM[41694] = 8'b10001011;
DRAM[41695] = 8'b10001010;
DRAM[41696] = 8'b10001100;
DRAM[41697] = 8'b10001001;
DRAM[41698] = 8'b10000110;
DRAM[41699] = 8'b10000101;
DRAM[41700] = 8'b10000101;
DRAM[41701] = 8'b10000101;
DRAM[41702] = 8'b10000101;
DRAM[41703] = 8'b10000100;
DRAM[41704] = 8'b10000000;
DRAM[41705] = 8'b10000000;
DRAM[41706] = 8'b1111110;
DRAM[41707] = 8'b1111101;
DRAM[41708] = 8'b1111100;
DRAM[41709] = 8'b1111100;
DRAM[41710] = 8'b1111100;
DRAM[41711] = 8'b1111101;
DRAM[41712] = 8'b1111100;
DRAM[41713] = 8'b1111101;
DRAM[41714] = 8'b1111111;
DRAM[41715] = 8'b10000010;
DRAM[41716] = 8'b10000011;
DRAM[41717] = 8'b10000011;
DRAM[41718] = 8'b10000010;
DRAM[41719] = 8'b10000010;
DRAM[41720] = 8'b10000110;
DRAM[41721] = 8'b10000100;
DRAM[41722] = 8'b10000001;
DRAM[41723] = 8'b10000001;
DRAM[41724] = 8'b10000001;
DRAM[41725] = 8'b10000001;
DRAM[41726] = 8'b10000000;
DRAM[41727] = 8'b1111111;
DRAM[41728] = 8'b10010111;
DRAM[41729] = 8'b10010111;
DRAM[41730] = 8'b10010111;
DRAM[41731] = 8'b10011000;
DRAM[41732] = 8'b10011000;
DRAM[41733] = 8'b10011001;
DRAM[41734] = 8'b10011001;
DRAM[41735] = 8'b10011001;
DRAM[41736] = 8'b10011100;
DRAM[41737] = 8'b10011101;
DRAM[41738] = 8'b10011110;
DRAM[41739] = 8'b10011111;
DRAM[41740] = 8'b10011111;
DRAM[41741] = 8'b10011111;
DRAM[41742] = 8'b10011111;
DRAM[41743] = 8'b10011111;
DRAM[41744] = 8'b10011110;
DRAM[41745] = 8'b10011110;
DRAM[41746] = 8'b10011111;
DRAM[41747] = 8'b10100000;
DRAM[41748] = 8'b10100001;
DRAM[41749] = 8'b10100010;
DRAM[41750] = 8'b10100010;
DRAM[41751] = 8'b10100011;
DRAM[41752] = 8'b10100011;
DRAM[41753] = 8'b10100100;
DRAM[41754] = 8'b10100100;
DRAM[41755] = 8'b10100100;
DRAM[41756] = 8'b10100100;
DRAM[41757] = 8'b10100101;
DRAM[41758] = 8'b10100101;
DRAM[41759] = 8'b10100101;
DRAM[41760] = 8'b10100100;
DRAM[41761] = 8'b10100011;
DRAM[41762] = 8'b10100001;
DRAM[41763] = 8'b10100001;
DRAM[41764] = 8'b10100100;
DRAM[41765] = 8'b10101000;
DRAM[41766] = 8'b10101011;
DRAM[41767] = 8'b10101101;
DRAM[41768] = 8'b10110011;
DRAM[41769] = 8'b11001000;
DRAM[41770] = 8'b11100010;
DRAM[41771] = 8'b11110101;
DRAM[41772] = 8'b11111101;
DRAM[41773] = 8'b11111111;
DRAM[41774] = 8'b11111110;
DRAM[41775] = 8'b11111010;
DRAM[41776] = 8'b11111110;
DRAM[41777] = 8'b11111110;
DRAM[41778] = 8'b11111110;
DRAM[41779] = 8'b11111110;
DRAM[41780] = 8'b11111110;
DRAM[41781] = 8'b11111110;
DRAM[41782] = 8'b11111110;
DRAM[41783] = 8'b11111110;
DRAM[41784] = 8'b11111111;
DRAM[41785] = 8'b11111110;
DRAM[41786] = 8'b11111101;
DRAM[41787] = 8'b11111101;
DRAM[41788] = 8'b11111101;
DRAM[41789] = 8'b11111011;
DRAM[41790] = 8'b11111000;
DRAM[41791] = 8'b11110101;
DRAM[41792] = 8'b11101111;
DRAM[41793] = 8'b11100111;
DRAM[41794] = 8'b11011100;
DRAM[41795] = 8'b11010101;
DRAM[41796] = 8'b11010001;
DRAM[41797] = 8'b11001110;
DRAM[41798] = 8'b11001011;
DRAM[41799] = 8'b11000111;
DRAM[41800] = 8'b10111110;
DRAM[41801] = 8'b10111100;
DRAM[41802] = 8'b10110011;
DRAM[41803] = 8'b10100111;
DRAM[41804] = 8'b10100001;
DRAM[41805] = 8'b10100010;
DRAM[41806] = 8'b10100100;
DRAM[41807] = 8'b10100100;
DRAM[41808] = 8'b10100000;
DRAM[41809] = 8'b10011101;
DRAM[41810] = 8'b10011001;
DRAM[41811] = 8'b10011000;
DRAM[41812] = 8'b10011001;
DRAM[41813] = 8'b10011010;
DRAM[41814] = 8'b10011010;
DRAM[41815] = 8'b10011001;
DRAM[41816] = 8'b10010010;
DRAM[41817] = 8'b10010110;
DRAM[41818] = 8'b10011111;
DRAM[41819] = 8'b10101011;
DRAM[41820] = 8'b10110011;
DRAM[41821] = 8'b10110100;
DRAM[41822] = 8'b10101100;
DRAM[41823] = 8'b10100101;
DRAM[41824] = 8'b10101000;
DRAM[41825] = 8'b10101001;
DRAM[41826] = 8'b10101011;
DRAM[41827] = 8'b10101101;
DRAM[41828] = 8'b10110001;
DRAM[41829] = 8'b10111000;
DRAM[41830] = 8'b11000000;
DRAM[41831] = 8'b11000110;
DRAM[41832] = 8'b11001000;
DRAM[41833] = 8'b11000111;
DRAM[41834] = 8'b11001000;
DRAM[41835] = 8'b11001100;
DRAM[41836] = 8'b11010001;
DRAM[41837] = 8'b11010100;
DRAM[41838] = 8'b11010011;
DRAM[41839] = 8'b11010000;
DRAM[41840] = 8'b11001111;
DRAM[41841] = 8'b11001101;
DRAM[41842] = 8'b11010100;
DRAM[41843] = 8'b11011000;
DRAM[41844] = 8'b11010110;
DRAM[41845] = 8'b11011001;
DRAM[41846] = 8'b11010011;
DRAM[41847] = 8'b11000011;
DRAM[41848] = 8'b10110111;
DRAM[41849] = 8'b11000001;
DRAM[41850] = 8'b10111101;
DRAM[41851] = 8'b10101100;
DRAM[41852] = 8'b10101010;
DRAM[41853] = 8'b10110111;
DRAM[41854] = 8'b10110111;
DRAM[41855] = 8'b10101011;
DRAM[41856] = 8'b10101000;
DRAM[41857] = 8'b10011111;
DRAM[41858] = 8'b10010101;
DRAM[41859] = 8'b10001000;
DRAM[41860] = 8'b1101110;
DRAM[41861] = 8'b1001011;
DRAM[41862] = 8'b101111;
DRAM[41863] = 8'b100100;
DRAM[41864] = 8'b100011;
DRAM[41865] = 8'b100001;
DRAM[41866] = 8'b100010;
DRAM[41867] = 8'b10110;
DRAM[41868] = 8'b11;
DRAM[41869] = 8'b0;
DRAM[41870] = 8'b101;
DRAM[41871] = 8'b0;
DRAM[41872] = 8'b0;
DRAM[41873] = 8'b0;
DRAM[41874] = 8'b0;
DRAM[41875] = 8'b0;
DRAM[41876] = 8'b0;
DRAM[41877] = 8'b0;
DRAM[41878] = 8'b0;
DRAM[41879] = 8'b0;
DRAM[41880] = 8'b0;
DRAM[41881] = 8'b0;
DRAM[41882] = 8'b0;
DRAM[41883] = 8'b0;
DRAM[41884] = 8'b0;
DRAM[41885] = 8'b11;
DRAM[41886] = 8'b1001;
DRAM[41887] = 8'b1110;
DRAM[41888] = 8'b11110;
DRAM[41889] = 8'b111001;
DRAM[41890] = 8'b1001100;
DRAM[41891] = 8'b1101010;
DRAM[41892] = 8'b10001010;
DRAM[41893] = 8'b10000011;
DRAM[41894] = 8'b10000000;
DRAM[41895] = 8'b10100001;
DRAM[41896] = 8'b10110011;
DRAM[41897] = 8'b10110011;
DRAM[41898] = 8'b10110110;
DRAM[41899] = 8'b10111100;
DRAM[41900] = 8'b11000000;
DRAM[41901] = 8'b11000101;
DRAM[41902] = 8'b11010000;
DRAM[41903] = 8'b11011100;
DRAM[41904] = 8'b11100011;
DRAM[41905] = 8'b11101001;
DRAM[41906] = 8'b11101001;
DRAM[41907] = 8'b11011111;
DRAM[41908] = 8'b11011001;
DRAM[41909] = 8'b11011011;
DRAM[41910] = 8'b11011100;
DRAM[41911] = 8'b11011010;
DRAM[41912] = 8'b11100001;
DRAM[41913] = 8'b11011100;
DRAM[41914] = 8'b11011101;
DRAM[41915] = 8'b11001100;
DRAM[41916] = 8'b11001001;
DRAM[41917] = 8'b11010010;
DRAM[41918] = 8'b11000101;
DRAM[41919] = 8'b11000010;
DRAM[41920] = 8'b11000101;
DRAM[41921] = 8'b11001010;
DRAM[41922] = 8'b11001110;
DRAM[41923] = 8'b11001111;
DRAM[41924] = 8'b11010001;
DRAM[41925] = 8'b11010000;
DRAM[41926] = 8'b11000101;
DRAM[41927] = 8'b10111000;
DRAM[41928] = 8'b11000000;
DRAM[41929] = 8'b10110101;
DRAM[41930] = 8'b10100111;
DRAM[41931] = 8'b10100000;
DRAM[41932] = 8'b10100101;
DRAM[41933] = 8'b10110011;
DRAM[41934] = 8'b11000001;
DRAM[41935] = 8'b11001001;
DRAM[41936] = 8'b10111010;
DRAM[41937] = 8'b10110010;
DRAM[41938] = 8'b10100111;
DRAM[41939] = 8'b10011101;
DRAM[41940] = 8'b10010111;
DRAM[41941] = 8'b10010100;
DRAM[41942] = 8'b10010011;
DRAM[41943] = 8'b10010010;
DRAM[41944] = 8'b10010110;
DRAM[41945] = 8'b10010101;
DRAM[41946] = 8'b10010100;
DRAM[41947] = 8'b10010010;
DRAM[41948] = 8'b10001111;
DRAM[41949] = 8'b10001101;
DRAM[41950] = 8'b10001011;
DRAM[41951] = 8'b10001001;
DRAM[41952] = 8'b10001011;
DRAM[41953] = 8'b10001000;
DRAM[41954] = 8'b10000101;
DRAM[41955] = 8'b10000100;
DRAM[41956] = 8'b10000100;
DRAM[41957] = 8'b10000100;
DRAM[41958] = 8'b10000011;
DRAM[41959] = 8'b10000010;
DRAM[41960] = 8'b1111111;
DRAM[41961] = 8'b1111111;
DRAM[41962] = 8'b1111110;
DRAM[41963] = 8'b1111101;
DRAM[41964] = 8'b1111100;
DRAM[41965] = 8'b1111100;
DRAM[41966] = 8'b1111100;
DRAM[41967] = 8'b1111101;
DRAM[41968] = 8'b1111101;
DRAM[41969] = 8'b1111110;
DRAM[41970] = 8'b1111111;
DRAM[41971] = 8'b10000001;
DRAM[41972] = 8'b10000011;
DRAM[41973] = 8'b10000011;
DRAM[41974] = 8'b10000011;
DRAM[41975] = 8'b10000011;
DRAM[41976] = 8'b10000111;
DRAM[41977] = 8'b10000101;
DRAM[41978] = 8'b10000011;
DRAM[41979] = 8'b10000010;
DRAM[41980] = 8'b10000010;
DRAM[41981] = 8'b10000010;
DRAM[41982] = 8'b10000001;
DRAM[41983] = 8'b1111111;
DRAM[41984] = 8'b10010111;
DRAM[41985] = 8'b10010111;
DRAM[41986] = 8'b10011000;
DRAM[41987] = 8'b10011000;
DRAM[41988] = 8'b10011000;
DRAM[41989] = 8'b10011000;
DRAM[41990] = 8'b10011001;
DRAM[41991] = 8'b10011001;
DRAM[41992] = 8'b10011011;
DRAM[41993] = 8'b10011100;
DRAM[41994] = 8'b10011101;
DRAM[41995] = 8'b10011110;
DRAM[41996] = 8'b10011111;
DRAM[41997] = 8'b10011111;
DRAM[41998] = 8'b10011111;
DRAM[41999] = 8'b10011110;
DRAM[42000] = 8'b10100000;
DRAM[42001] = 8'b10100000;
DRAM[42002] = 8'b10100001;
DRAM[42003] = 8'b10100001;
DRAM[42004] = 8'b10100010;
DRAM[42005] = 8'b10100011;
DRAM[42006] = 8'b10100011;
DRAM[42007] = 8'b10100011;
DRAM[42008] = 8'b10100010;
DRAM[42009] = 8'b10100011;
DRAM[42010] = 8'b10100011;
DRAM[42011] = 8'b10100100;
DRAM[42012] = 8'b10100100;
DRAM[42013] = 8'b10100101;
DRAM[42014] = 8'b10100101;
DRAM[42015] = 8'b10100101;
DRAM[42016] = 8'b10100011;
DRAM[42017] = 8'b10100100;
DRAM[42018] = 8'b10100101;
DRAM[42019] = 8'b10100111;
DRAM[42020] = 8'b10101001;
DRAM[42021] = 8'b10101101;
DRAM[42022] = 8'b10110010;
DRAM[42023] = 8'b10110101;
DRAM[42024] = 8'b10111110;
DRAM[42025] = 8'b11011010;
DRAM[42026] = 8'b11110110;
DRAM[42027] = 8'b11111111;
DRAM[42028] = 8'b11111110;
DRAM[42029] = 8'b11111101;
DRAM[42030] = 8'b11111110;
DRAM[42031] = 8'b11111110;
DRAM[42032] = 8'b11111110;
DRAM[42033] = 8'b11111110;
DRAM[42034] = 8'b11111110;
DRAM[42035] = 8'b11111110;
DRAM[42036] = 8'b11111110;
DRAM[42037] = 8'b11111110;
DRAM[42038] = 8'b11111110;
DRAM[42039] = 8'b11111110;
DRAM[42040] = 8'b11111111;
DRAM[42041] = 8'b11111110;
DRAM[42042] = 8'b11111101;
DRAM[42043] = 8'b11111100;
DRAM[42044] = 8'b11111100;
DRAM[42045] = 8'b11111010;
DRAM[42046] = 8'b11110110;
DRAM[42047] = 8'b11110011;
DRAM[42048] = 8'b11101100;
DRAM[42049] = 8'b11100100;
DRAM[42050] = 8'b11011010;
DRAM[42051] = 8'b11010011;
DRAM[42052] = 8'b11001111;
DRAM[42053] = 8'b11001100;
DRAM[42054] = 8'b11001001;
DRAM[42055] = 8'b11000110;
DRAM[42056] = 8'b11000011;
DRAM[42057] = 8'b10111110;
DRAM[42058] = 8'b10110101;
DRAM[42059] = 8'b10101101;
DRAM[42060] = 8'b10101110;
DRAM[42061] = 8'b10110010;
DRAM[42062] = 8'b10110001;
DRAM[42063] = 8'b10101100;
DRAM[42064] = 8'b10100001;
DRAM[42065] = 8'b10011101;
DRAM[42066] = 8'b10010111;
DRAM[42067] = 8'b10010011;
DRAM[42068] = 8'b10010010;
DRAM[42069] = 8'b10010001;
DRAM[42070] = 8'b10010001;
DRAM[42071] = 8'b10010000;
DRAM[42072] = 8'b10010101;
DRAM[42073] = 8'b10010101;
DRAM[42074] = 8'b10010101;
DRAM[42075] = 8'b10010111;
DRAM[42076] = 8'b10011100;
DRAM[42077] = 8'b10100100;
DRAM[42078] = 8'b10101101;
DRAM[42079] = 8'b10110010;
DRAM[42080] = 8'b10101101;
DRAM[42081] = 8'b10101101;
DRAM[42082] = 8'b10101111;
DRAM[42083] = 8'b10110000;
DRAM[42084] = 8'b10110100;
DRAM[42085] = 8'b10111011;
DRAM[42086] = 8'b11000011;
DRAM[42087] = 8'b11001001;
DRAM[42088] = 8'b11010011;
DRAM[42089] = 8'b11010000;
DRAM[42090] = 8'b11001101;
DRAM[42091] = 8'b11001110;
DRAM[42092] = 8'b11010000;
DRAM[42093] = 8'b11010000;
DRAM[42094] = 8'b11001101;
DRAM[42095] = 8'b11001010;
DRAM[42096] = 8'b11001101;
DRAM[42097] = 8'b11010010;
DRAM[42098] = 8'b11011100;
DRAM[42099] = 8'b11011000;
DRAM[42100] = 8'b11001001;
DRAM[42101] = 8'b11001001;
DRAM[42102] = 8'b11001111;
DRAM[42103] = 8'b11001011;
DRAM[42104] = 8'b11001001;
DRAM[42105] = 8'b11010000;
DRAM[42106] = 8'b11001010;
DRAM[42107] = 8'b10111011;
DRAM[42108] = 8'b10111001;
DRAM[42109] = 8'b10111110;
DRAM[42110] = 8'b10110000;
DRAM[42111] = 8'b10011001;
DRAM[42112] = 8'b10010110;
DRAM[42113] = 8'b10010100;
DRAM[42114] = 8'b10010011;
DRAM[42115] = 8'b10001101;
DRAM[42116] = 8'b1111011;
DRAM[42117] = 8'b1011010;
DRAM[42118] = 8'b110101;
DRAM[42119] = 8'b11101;
DRAM[42120] = 8'b11010;
DRAM[42121] = 8'b10100;
DRAM[42122] = 8'b10010;
DRAM[42123] = 8'b1000;
DRAM[42124] = 8'b0;
DRAM[42125] = 8'b0;
DRAM[42126] = 8'b10;
DRAM[42127] = 8'b0;
DRAM[42128] = 8'b0;
DRAM[42129] = 8'b0;
DRAM[42130] = 8'b0;
DRAM[42131] = 8'b0;
DRAM[42132] = 8'b0;
DRAM[42133] = 8'b0;
DRAM[42134] = 8'b0;
DRAM[42135] = 8'b0;
DRAM[42136] = 8'b1;
DRAM[42137] = 8'b10;
DRAM[42138] = 8'b11;
DRAM[42139] = 8'b11;
DRAM[42140] = 8'b11;
DRAM[42141] = 8'b101;
DRAM[42142] = 8'b111;
DRAM[42143] = 8'b1010;
DRAM[42144] = 8'b11001;
DRAM[42145] = 8'b111001;
DRAM[42146] = 8'b1001101;
DRAM[42147] = 8'b1100100;
DRAM[42148] = 8'b1111101;
DRAM[42149] = 8'b1110110;
DRAM[42150] = 8'b1111001;
DRAM[42151] = 8'b10011110;
DRAM[42152] = 8'b10110001;
DRAM[42153] = 8'b10101111;
DRAM[42154] = 8'b10101111;
DRAM[42155] = 8'b10110001;
DRAM[42156] = 8'b10110010;
DRAM[42157] = 8'b10110110;
DRAM[42158] = 8'b11000010;
DRAM[42159] = 8'b11001101;
DRAM[42160] = 8'b11011110;
DRAM[42161] = 8'b11101011;
DRAM[42162] = 8'b11101110;
DRAM[42163] = 8'b11011111;
DRAM[42164] = 8'b11010010;
DRAM[42165] = 8'b11010001;
DRAM[42166] = 8'b11010101;
DRAM[42167] = 8'b11010101;
DRAM[42168] = 8'b11010011;
DRAM[42169] = 8'b11001101;
DRAM[42170] = 8'b11001101;
DRAM[42171] = 8'b10111100;
DRAM[42172] = 8'b10111011;
DRAM[42173] = 8'b11001000;
DRAM[42174] = 8'b11000000;
DRAM[42175] = 8'b10111111;
DRAM[42176] = 8'b11001100;
DRAM[42177] = 8'b11010010;
DRAM[42178] = 8'b11010100;
DRAM[42179] = 8'b11001101;
DRAM[42180] = 8'b11000110;
DRAM[42181] = 8'b11000110;
DRAM[42182] = 8'b11001100;
DRAM[42183] = 8'b11010001;
DRAM[42184] = 8'b10111101;
DRAM[42185] = 8'b10110100;
DRAM[42186] = 8'b10101011;
DRAM[42187] = 8'b10101001;
DRAM[42188] = 8'b10101011;
DRAM[42189] = 8'b10101010;
DRAM[42190] = 8'b10100100;
DRAM[42191] = 8'b10011110;
DRAM[42192] = 8'b10110010;
DRAM[42193] = 8'b10110011;
DRAM[42194] = 8'b10110100;
DRAM[42195] = 8'b10110011;
DRAM[42196] = 8'b10101111;
DRAM[42197] = 8'b10100101;
DRAM[42198] = 8'b10011010;
DRAM[42199] = 8'b10010001;
DRAM[42200] = 8'b10010010;
DRAM[42201] = 8'b10010010;
DRAM[42202] = 8'b10010011;
DRAM[42203] = 8'b10010011;
DRAM[42204] = 8'b10010011;
DRAM[42205] = 8'b10010001;
DRAM[42206] = 8'b10010000;
DRAM[42207] = 8'b10001111;
DRAM[42208] = 8'b10001000;
DRAM[42209] = 8'b10000101;
DRAM[42210] = 8'b10000011;
DRAM[42211] = 8'b10000010;
DRAM[42212] = 8'b10000011;
DRAM[42213] = 8'b10000010;
DRAM[42214] = 8'b10000001;
DRAM[42215] = 8'b1111111;
DRAM[42216] = 8'b1111110;
DRAM[42217] = 8'b1111110;
DRAM[42218] = 8'b1111101;
DRAM[42219] = 8'b1111100;
DRAM[42220] = 8'b1111100;
DRAM[42221] = 8'b1111100;
DRAM[42222] = 8'b1111100;
DRAM[42223] = 8'b1111101;
DRAM[42224] = 8'b1111110;
DRAM[42225] = 8'b1111110;
DRAM[42226] = 8'b10000000;
DRAM[42227] = 8'b10000001;
DRAM[42228] = 8'b10000010;
DRAM[42229] = 8'b10000011;
DRAM[42230] = 8'b10000100;
DRAM[42231] = 8'b10000100;
DRAM[42232] = 8'b10000111;
DRAM[42233] = 8'b10000101;
DRAM[42234] = 8'b10000011;
DRAM[42235] = 8'b10000011;
DRAM[42236] = 8'b10000100;
DRAM[42237] = 8'b10000100;
DRAM[42238] = 8'b10000010;
DRAM[42239] = 8'b10000000;
DRAM[42240] = 8'b10011000;
DRAM[42241] = 8'b10011000;
DRAM[42242] = 8'b10011000;
DRAM[42243] = 8'b10011000;
DRAM[42244] = 8'b10011000;
DRAM[42245] = 8'b10011000;
DRAM[42246] = 8'b10011000;
DRAM[42247] = 8'b10011000;
DRAM[42248] = 8'b10011010;
DRAM[42249] = 8'b10011011;
DRAM[42250] = 8'b10011100;
DRAM[42251] = 8'b10011110;
DRAM[42252] = 8'b10011111;
DRAM[42253] = 8'b10011111;
DRAM[42254] = 8'b10011111;
DRAM[42255] = 8'b10011111;
DRAM[42256] = 8'b10100001;
DRAM[42257] = 8'b10100001;
DRAM[42258] = 8'b10100010;
DRAM[42259] = 8'b10100010;
DRAM[42260] = 8'b10100010;
DRAM[42261] = 8'b10100011;
DRAM[42262] = 8'b10100011;
DRAM[42263] = 8'b10100011;
DRAM[42264] = 8'b10100010;
DRAM[42265] = 8'b10100010;
DRAM[42266] = 8'b10100010;
DRAM[42267] = 8'b10100011;
DRAM[42268] = 8'b10100100;
DRAM[42269] = 8'b10100100;
DRAM[42270] = 8'b10100101;
DRAM[42271] = 8'b10100101;
DRAM[42272] = 8'b10100000;
DRAM[42273] = 8'b10100100;
DRAM[42274] = 8'b10100111;
DRAM[42275] = 8'b10100110;
DRAM[42276] = 8'b10100101;
DRAM[42277] = 8'b10101000;
DRAM[42278] = 8'b10110001;
DRAM[42279] = 8'b10111001;
DRAM[42280] = 8'b11010000;
DRAM[42281] = 8'b11101001;
DRAM[42282] = 8'b11111110;
DRAM[42283] = 8'b11111111;
DRAM[42284] = 8'b11111011;
DRAM[42285] = 8'b11111100;
DRAM[42286] = 8'b11111111;
DRAM[42287] = 8'b11111111;
DRAM[42288] = 8'b11111110;
DRAM[42289] = 8'b11111110;
DRAM[42290] = 8'b11111110;
DRAM[42291] = 8'b11111110;
DRAM[42292] = 8'b11111110;
DRAM[42293] = 8'b11111110;
DRAM[42294] = 8'b11111110;
DRAM[42295] = 8'b11111110;
DRAM[42296] = 8'b11111111;
DRAM[42297] = 8'b11111110;
DRAM[42298] = 8'b11111100;
DRAM[42299] = 8'b11111100;
DRAM[42300] = 8'b11111011;
DRAM[42301] = 8'b11111001;
DRAM[42302] = 8'b11110100;
DRAM[42303] = 8'b11110001;
DRAM[42304] = 8'b11101010;
DRAM[42305] = 8'b11100011;
DRAM[42306] = 8'b11011001;
DRAM[42307] = 8'b11010010;
DRAM[42308] = 8'b11001111;
DRAM[42309] = 8'b11001011;
DRAM[42310] = 8'b11000111;
DRAM[42311] = 8'b11000011;
DRAM[42312] = 8'b11000010;
DRAM[42313] = 8'b11000000;
DRAM[42314] = 8'b10111100;
DRAM[42315] = 8'b10111001;
DRAM[42316] = 8'b10111010;
DRAM[42317] = 8'b10111001;
DRAM[42318] = 8'b10101111;
DRAM[42319] = 8'b10100011;
DRAM[42320] = 8'b10011011;
DRAM[42321] = 8'b10010111;
DRAM[42322] = 8'b10010001;
DRAM[42323] = 8'b10001110;
DRAM[42324] = 8'b10001101;
DRAM[42325] = 8'b10001101;
DRAM[42326] = 8'b10001101;
DRAM[42327] = 8'b10001101;
DRAM[42328] = 8'b10010010;
DRAM[42329] = 8'b10010110;
DRAM[42330] = 8'b10011001;
DRAM[42331] = 8'b10011001;
DRAM[42332] = 8'b10011001;
DRAM[42333] = 8'b10011101;
DRAM[42334] = 8'b10100110;
DRAM[42335] = 8'b10101101;
DRAM[42336] = 8'b10100101;
DRAM[42337] = 8'b10101001;
DRAM[42338] = 8'b10110000;
DRAM[42339] = 8'b10110101;
DRAM[42340] = 8'b10111000;
DRAM[42341] = 8'b10111011;
DRAM[42342] = 8'b10111101;
DRAM[42343] = 8'b10111111;
DRAM[42344] = 8'b11001101;
DRAM[42345] = 8'b11001101;
DRAM[42346] = 8'b11001101;
DRAM[42347] = 8'b11001111;
DRAM[42348] = 8'b11010000;
DRAM[42349] = 8'b11010001;
DRAM[42350] = 8'b11010000;
DRAM[42351] = 8'b11001110;
DRAM[42352] = 8'b11010001;
DRAM[42353] = 8'b11011000;
DRAM[42354] = 8'b11100001;
DRAM[42355] = 8'b11010110;
DRAM[42356] = 8'b10111110;
DRAM[42357] = 8'b10111001;
DRAM[42358] = 8'b11000010;
DRAM[42359] = 8'b11000100;
DRAM[42360] = 8'b11000110;
DRAM[42361] = 8'b11000111;
DRAM[42362] = 8'b11000000;
DRAM[42363] = 8'b10110111;
DRAM[42364] = 8'b10110111;
DRAM[42365] = 8'b10110111;
DRAM[42366] = 8'b10100110;
DRAM[42367] = 8'b10001110;
DRAM[42368] = 8'b10000011;
DRAM[42369] = 8'b10001100;
DRAM[42370] = 8'b10010001;
DRAM[42371] = 8'b10001000;
DRAM[42372] = 8'b1110011;
DRAM[42373] = 8'b1010110;
DRAM[42374] = 8'b111010;
DRAM[42375] = 8'b100111;
DRAM[42376] = 8'b11011;
DRAM[42377] = 8'b1100;
DRAM[42378] = 8'b101;
DRAM[42379] = 8'b11;
DRAM[42380] = 8'b0;
DRAM[42381] = 8'b1;
DRAM[42382] = 8'b100;
DRAM[42383] = 8'b0;
DRAM[42384] = 8'b0;
DRAM[42385] = 8'b0;
DRAM[42386] = 8'b0;
DRAM[42387] = 8'b0;
DRAM[42388] = 8'b0;
DRAM[42389] = 8'b0;
DRAM[42390] = 8'b0;
DRAM[42391] = 8'b0;
DRAM[42392] = 8'b0;
DRAM[42393] = 8'b1;
DRAM[42394] = 8'b1;
DRAM[42395] = 8'b10;
DRAM[42396] = 8'b11;
DRAM[42397] = 8'b100;
DRAM[42398] = 8'b100;
DRAM[42399] = 8'b101;
DRAM[42400] = 8'b1111;
DRAM[42401] = 8'b110001;
DRAM[42402] = 8'b1001101;
DRAM[42403] = 8'b1100100;
DRAM[42404] = 8'b1111000;
DRAM[42405] = 8'b1111010;
DRAM[42406] = 8'b10000011;
DRAM[42407] = 8'b10011110;
DRAM[42408] = 8'b10100100;
DRAM[42409] = 8'b10100100;
DRAM[42410] = 8'b10100111;
DRAM[42411] = 8'b10101110;
DRAM[42412] = 8'b10110011;
DRAM[42413] = 8'b10111010;
DRAM[42414] = 8'b11000110;
DRAM[42415] = 8'b11010011;
DRAM[42416] = 8'b11010111;
DRAM[42417] = 8'b11101001;
DRAM[42418] = 8'b11110000;
DRAM[42419] = 8'b11011111;
DRAM[42420] = 8'b11001111;
DRAM[42421] = 8'b11001111;
DRAM[42422] = 8'b11010011;
DRAM[42423] = 8'b11010011;
DRAM[42424] = 8'b11011011;
DRAM[42425] = 8'b11011110;
DRAM[42426] = 8'b11100100;
DRAM[42427] = 8'b11001010;
DRAM[42428] = 8'b10111001;
DRAM[42429] = 8'b10111111;
DRAM[42430] = 8'b10111111;
DRAM[42431] = 8'b11001010;
DRAM[42432] = 8'b11001001;
DRAM[42433] = 8'b11001100;
DRAM[42434] = 8'b11001111;
DRAM[42435] = 8'b11010001;
DRAM[42436] = 8'b11010010;
DRAM[42437] = 8'b11010000;
DRAM[42438] = 8'b11001100;
DRAM[42439] = 8'b11001001;
DRAM[42440] = 8'b11010110;
DRAM[42441] = 8'b11001000;
DRAM[42442] = 8'b10110110;
DRAM[42443] = 8'b10100111;
DRAM[42444] = 8'b10100000;
DRAM[42445] = 8'b10011111;
DRAM[42446] = 8'b10011110;
DRAM[42447] = 8'b10011101;
DRAM[42448] = 8'b10010111;
DRAM[42449] = 8'b10011010;
DRAM[42450] = 8'b10100000;
DRAM[42451] = 8'b10100111;
DRAM[42452] = 8'b10101100;
DRAM[42453] = 8'b10101110;
DRAM[42454] = 8'b10101100;
DRAM[42455] = 8'b10101010;
DRAM[42456] = 8'b10011010;
DRAM[42457] = 8'b10011010;
DRAM[42458] = 8'b10011001;
DRAM[42459] = 8'b10010111;
DRAM[42460] = 8'b10010100;
DRAM[42461] = 8'b10010000;
DRAM[42462] = 8'b10001100;
DRAM[42463] = 8'b10001010;
DRAM[42464] = 8'b10000110;
DRAM[42465] = 8'b10000100;
DRAM[42466] = 8'b10000010;
DRAM[42467] = 8'b10000010;
DRAM[42468] = 8'b10000010;
DRAM[42469] = 8'b10000001;
DRAM[42470] = 8'b1111111;
DRAM[42471] = 8'b1111101;
DRAM[42472] = 8'b1111101;
DRAM[42473] = 8'b1111101;
DRAM[42474] = 8'b1111100;
DRAM[42475] = 8'b1111100;
DRAM[42476] = 8'b1111100;
DRAM[42477] = 8'b1111100;
DRAM[42478] = 8'b1111101;
DRAM[42479] = 8'b1111101;
DRAM[42480] = 8'b1111111;
DRAM[42481] = 8'b1111111;
DRAM[42482] = 8'b10000000;
DRAM[42483] = 8'b10000001;
DRAM[42484] = 8'b10000010;
DRAM[42485] = 8'b10000011;
DRAM[42486] = 8'b10000100;
DRAM[42487] = 8'b10000101;
DRAM[42488] = 8'b10000101;
DRAM[42489] = 8'b10000100;
DRAM[42490] = 8'b10000100;
DRAM[42491] = 8'b10000100;
DRAM[42492] = 8'b10000110;
DRAM[42493] = 8'b10000101;
DRAM[42494] = 8'b10000011;
DRAM[42495] = 8'b10000001;
DRAM[42496] = 8'b10011000;
DRAM[42497] = 8'b10011000;
DRAM[42498] = 8'b10011000;
DRAM[42499] = 8'b10011000;
DRAM[42500] = 8'b10011000;
DRAM[42501] = 8'b10011000;
DRAM[42502] = 8'b10011000;
DRAM[42503] = 8'b10011000;
DRAM[42504] = 8'b10011001;
DRAM[42505] = 8'b10011010;
DRAM[42506] = 8'b10011011;
DRAM[42507] = 8'b10011101;
DRAM[42508] = 8'b10011111;
DRAM[42509] = 8'b10100000;
DRAM[42510] = 8'b10100000;
DRAM[42511] = 8'b10100000;
DRAM[42512] = 8'b10100000;
DRAM[42513] = 8'b10100001;
DRAM[42514] = 8'b10100001;
DRAM[42515] = 8'b10100001;
DRAM[42516] = 8'b10100001;
DRAM[42517] = 8'b10100010;
DRAM[42518] = 8'b10100010;
DRAM[42519] = 8'b10100010;
DRAM[42520] = 8'b10100001;
DRAM[42521] = 8'b10100001;
DRAM[42522] = 8'b10100010;
DRAM[42523] = 8'b10100011;
DRAM[42524] = 8'b10100100;
DRAM[42525] = 8'b10100100;
DRAM[42526] = 8'b10100101;
DRAM[42527] = 8'b10100101;
DRAM[42528] = 8'b10100000;
DRAM[42529] = 8'b10100110;
DRAM[42530] = 8'b10101000;
DRAM[42531] = 8'b10100101;
DRAM[42532] = 8'b10100001;
DRAM[42533] = 8'b10100110;
DRAM[42534] = 8'b10110111;
DRAM[42535] = 8'b11000110;
DRAM[42536] = 8'b11100100;
DRAM[42537] = 8'b11110100;
DRAM[42538] = 8'b11111110;
DRAM[42539] = 8'b11111100;
DRAM[42540] = 8'b11111011;
DRAM[42541] = 8'b11111111;
DRAM[42542] = 8'b11111111;
DRAM[42543] = 8'b11111100;
DRAM[42544] = 8'b11111110;
DRAM[42545] = 8'b11111110;
DRAM[42546] = 8'b11111110;
DRAM[42547] = 8'b11111110;
DRAM[42548] = 8'b11111110;
DRAM[42549] = 8'b11111110;
DRAM[42550] = 8'b11111110;
DRAM[42551] = 8'b11111110;
DRAM[42552] = 8'b11111111;
DRAM[42553] = 8'b11111110;
DRAM[42554] = 8'b11111100;
DRAM[42555] = 8'b11111011;
DRAM[42556] = 8'b11111010;
DRAM[42557] = 8'b11111000;
DRAM[42558] = 8'b11110011;
DRAM[42559] = 8'b11110000;
DRAM[42560] = 8'b11101010;
DRAM[42561] = 8'b11100100;
DRAM[42562] = 8'b11011011;
DRAM[42563] = 8'b11010100;
DRAM[42564] = 8'b11010000;
DRAM[42565] = 8'b11001100;
DRAM[42566] = 8'b11000110;
DRAM[42567] = 8'b11000001;
DRAM[42568] = 8'b10111110;
DRAM[42569] = 8'b11000000;
DRAM[42570] = 8'b10111110;
DRAM[42571] = 8'b10111010;
DRAM[42572] = 8'b10110110;
DRAM[42573] = 8'b10110000;
DRAM[42574] = 8'b10100101;
DRAM[42575] = 8'b10011010;
DRAM[42576] = 8'b10011011;
DRAM[42577] = 8'b10010111;
DRAM[42578] = 8'b10010010;
DRAM[42579] = 8'b10001111;
DRAM[42580] = 8'b10001111;
DRAM[42581] = 8'b10001111;
DRAM[42582] = 8'b10001111;
DRAM[42583] = 8'b10001110;
DRAM[42584] = 8'b10001011;
DRAM[42585] = 8'b10010011;
DRAM[42586] = 8'b10011100;
DRAM[42587] = 8'b10100001;
DRAM[42588] = 8'b10100001;
DRAM[42589] = 8'b10100000;
DRAM[42590] = 8'b10100000;
DRAM[42591] = 8'b10100010;
DRAM[42592] = 8'b10100011;
DRAM[42593] = 8'b10101000;
DRAM[42594] = 8'b10110000;
DRAM[42595] = 8'b10110101;
DRAM[42596] = 8'b10111001;
DRAM[42597] = 8'b10111011;
DRAM[42598] = 8'b10111101;
DRAM[42599] = 8'b10111110;
DRAM[42600] = 8'b11000010;
DRAM[42601] = 8'b11000110;
DRAM[42602] = 8'b11001010;
DRAM[42603] = 8'b11001110;
DRAM[42604] = 8'b11010000;
DRAM[42605] = 8'b11010010;
DRAM[42606] = 8'b11010100;
DRAM[42607] = 8'b11010101;
DRAM[42608] = 8'b11010100;
DRAM[42609] = 8'b11010110;
DRAM[42610] = 8'b11011010;
DRAM[42611] = 8'b11001111;
DRAM[42612] = 8'b10111001;
DRAM[42613] = 8'b10110100;
DRAM[42614] = 8'b10110111;
DRAM[42615] = 8'b10110011;
DRAM[42616] = 8'b10110010;
DRAM[42617] = 8'b10101110;
DRAM[42618] = 8'b10101000;
DRAM[42619] = 8'b10100101;
DRAM[42620] = 8'b10100111;
DRAM[42621] = 8'b10101001;
DRAM[42622] = 8'b10100001;
DRAM[42623] = 8'b10010101;
DRAM[42624] = 8'b10000111;
DRAM[42625] = 8'b10001001;
DRAM[42626] = 8'b10000100;
DRAM[42627] = 8'b1110101;
DRAM[42628] = 8'b1100100;
DRAM[42629] = 8'b1010100;
DRAM[42630] = 8'b1000001;
DRAM[42631] = 8'b110000;
DRAM[42632] = 8'b100000;
DRAM[42633] = 8'b1010;
DRAM[42634] = 8'b10;
DRAM[42635] = 8'b110;
DRAM[42636] = 8'b11;
DRAM[42637] = 8'b11;
DRAM[42638] = 8'b101;
DRAM[42639] = 8'b1;
DRAM[42640] = 8'b0;
DRAM[42641] = 8'b0;
DRAM[42642] = 8'b0;
DRAM[42643] = 8'b0;
DRAM[42644] = 8'b0;
DRAM[42645] = 8'b0;
DRAM[42646] = 8'b0;
DRAM[42647] = 8'b0;
DRAM[42648] = 8'b0;
DRAM[42649] = 8'b0;
DRAM[42650] = 8'b0;
DRAM[42651] = 8'b0;
DRAM[42652] = 8'b1;
DRAM[42653] = 8'b1;
DRAM[42654] = 8'b0;
DRAM[42655] = 8'b0;
DRAM[42656] = 8'b10001;
DRAM[42657] = 8'b101110;
DRAM[42658] = 8'b1001101;
DRAM[42659] = 8'b1011111;
DRAM[42660] = 8'b1101100;
DRAM[42661] = 8'b1111011;
DRAM[42662] = 8'b10001101;
DRAM[42663] = 8'b10011010;
DRAM[42664] = 8'b10011100;
DRAM[42665] = 8'b10011110;
DRAM[42666] = 8'b10100110;
DRAM[42667] = 8'b10110001;
DRAM[42668] = 8'b10111001;
DRAM[42669] = 8'b11000001;
DRAM[42670] = 8'b11001101;
DRAM[42671] = 8'b11011001;
DRAM[42672] = 8'b11010101;
DRAM[42673] = 8'b11101000;
DRAM[42674] = 8'b11101110;
DRAM[42675] = 8'b11011111;
DRAM[42676] = 8'b11010010;
DRAM[42677] = 8'b11010011;
DRAM[42678] = 8'b11010100;
DRAM[42679] = 8'b11010000;
DRAM[42680] = 8'b11010101;
DRAM[42681] = 8'b11011011;
DRAM[42682] = 8'b11100010;
DRAM[42683] = 8'b11000111;
DRAM[42684] = 8'b10110010;
DRAM[42685] = 8'b10110100;
DRAM[42686] = 8'b10110011;
DRAM[42687] = 8'b10111111;
DRAM[42688] = 8'b11011111;
DRAM[42689] = 8'b11010000;
DRAM[42690] = 8'b11000000;
DRAM[42691] = 8'b10111100;
DRAM[42692] = 8'b11000001;
DRAM[42693] = 8'b11001000;
DRAM[42694] = 8'b11001001;
DRAM[42695] = 8'b11001000;
DRAM[42696] = 8'b11001000;
DRAM[42697] = 8'b11000111;
DRAM[42698] = 8'b11000001;
DRAM[42699] = 8'b10110100;
DRAM[42700] = 8'b10100110;
DRAM[42701] = 8'b10100000;
DRAM[42702] = 8'b10100011;
DRAM[42703] = 8'b10101000;
DRAM[42704] = 8'b10100011;
DRAM[42705] = 8'b10011110;
DRAM[42706] = 8'b10011000;
DRAM[42707] = 8'b10010101;
DRAM[42708] = 8'b10010110;
DRAM[42709] = 8'b10011000;
DRAM[42710] = 8'b10011010;
DRAM[42711] = 8'b10011100;
DRAM[42712] = 8'b10011110;
DRAM[42713] = 8'b10011110;
DRAM[42714] = 8'b10011101;
DRAM[42715] = 8'b10011010;
DRAM[42716] = 8'b10010110;
DRAM[42717] = 8'b10010001;
DRAM[42718] = 8'b10001100;
DRAM[42719] = 8'b10001010;
DRAM[42720] = 8'b10000110;
DRAM[42721] = 8'b10000100;
DRAM[42722] = 8'b10000011;
DRAM[42723] = 8'b10000010;
DRAM[42724] = 8'b10000011;
DRAM[42725] = 8'b10000010;
DRAM[42726] = 8'b1111111;
DRAM[42727] = 8'b1111101;
DRAM[42728] = 8'b1111101;
DRAM[42729] = 8'b1111100;
DRAM[42730] = 8'b1111100;
DRAM[42731] = 8'b1111011;
DRAM[42732] = 8'b1111011;
DRAM[42733] = 8'b1111100;
DRAM[42734] = 8'b1111101;
DRAM[42735] = 8'b1111101;
DRAM[42736] = 8'b1111111;
DRAM[42737] = 8'b1111111;
DRAM[42738] = 8'b10000000;
DRAM[42739] = 8'b10000001;
DRAM[42740] = 8'b10000010;
DRAM[42741] = 8'b10000011;
DRAM[42742] = 8'b10000101;
DRAM[42743] = 8'b10000110;
DRAM[42744] = 8'b10000100;
DRAM[42745] = 8'b10000011;
DRAM[42746] = 8'b10000011;
DRAM[42747] = 8'b10000101;
DRAM[42748] = 8'b10000111;
DRAM[42749] = 8'b10000111;
DRAM[42750] = 8'b10000101;
DRAM[42751] = 8'b10000011;
DRAM[42752] = 8'b10011000;
DRAM[42753] = 8'b10011000;
DRAM[42754] = 8'b10011000;
DRAM[42755] = 8'b10011000;
DRAM[42756] = 8'b10011000;
DRAM[42757] = 8'b10011000;
DRAM[42758] = 8'b10011000;
DRAM[42759] = 8'b10011000;
DRAM[42760] = 8'b10010111;
DRAM[42761] = 8'b10011001;
DRAM[42762] = 8'b10011011;
DRAM[42763] = 8'b10011101;
DRAM[42764] = 8'b10011111;
DRAM[42765] = 8'b10100000;
DRAM[42766] = 8'b10100001;
DRAM[42767] = 8'b10100001;
DRAM[42768] = 8'b10011111;
DRAM[42769] = 8'b10011111;
DRAM[42770] = 8'b10100000;
DRAM[42771] = 8'b10100000;
DRAM[42772] = 8'b10100000;
DRAM[42773] = 8'b10100000;
DRAM[42774] = 8'b10100001;
DRAM[42775] = 8'b10100001;
DRAM[42776] = 8'b10100000;
DRAM[42777] = 8'b10100001;
DRAM[42778] = 8'b10100010;
DRAM[42779] = 8'b10100010;
DRAM[42780] = 8'b10100011;
DRAM[42781] = 8'b10100100;
DRAM[42782] = 8'b10100101;
DRAM[42783] = 8'b10100101;
DRAM[42784] = 8'b10100101;
DRAM[42785] = 8'b10101100;
DRAM[42786] = 8'b10101110;
DRAM[42787] = 8'b10101001;
DRAM[42788] = 8'b10100101;
DRAM[42789] = 8'b10101111;
DRAM[42790] = 8'b11000111;
DRAM[42791] = 8'b11011100;
DRAM[42792] = 8'b11110001;
DRAM[42793] = 8'b11111001;
DRAM[42794] = 8'b11111011;
DRAM[42795] = 8'b11111000;
DRAM[42796] = 8'b11111101;
DRAM[42797] = 8'b11111111;
DRAM[42798] = 8'b11111111;
DRAM[42799] = 8'b11110111;
DRAM[42800] = 8'b11111110;
DRAM[42801] = 8'b11111110;
DRAM[42802] = 8'b11111110;
DRAM[42803] = 8'b11111110;
DRAM[42804] = 8'b11111110;
DRAM[42805] = 8'b11111110;
DRAM[42806] = 8'b11111110;
DRAM[42807] = 8'b11111110;
DRAM[42808] = 8'b11111111;
DRAM[42809] = 8'b11111110;
DRAM[42810] = 8'b11111100;
DRAM[42811] = 8'b11111011;
DRAM[42812] = 8'b11111010;
DRAM[42813] = 8'b11110111;
DRAM[42814] = 8'b11110011;
DRAM[42815] = 8'b11101111;
DRAM[42816] = 8'b11101011;
DRAM[42817] = 8'b11100101;
DRAM[42818] = 8'b11011101;
DRAM[42819] = 8'b11010110;
DRAM[42820] = 8'b11010010;
DRAM[42821] = 8'b11001101;
DRAM[42822] = 8'b11000110;
DRAM[42823] = 8'b11000000;
DRAM[42824] = 8'b11000000;
DRAM[42825] = 8'b11000011;
DRAM[42826] = 8'b11000000;
DRAM[42827] = 8'b10110110;
DRAM[42828] = 8'b10101101;
DRAM[42829] = 8'b10101000;
DRAM[42830] = 8'b10100100;
DRAM[42831] = 8'b10011111;
DRAM[42832] = 8'b10100000;
DRAM[42833] = 8'b10011100;
DRAM[42834] = 8'b10011000;
DRAM[42835] = 8'b10010100;
DRAM[42836] = 8'b10010011;
DRAM[42837] = 8'b10010011;
DRAM[42838] = 8'b10010010;
DRAM[42839] = 8'b10010000;
DRAM[42840] = 8'b10010000;
DRAM[42841] = 8'b10010010;
DRAM[42842] = 8'b10010100;
DRAM[42843] = 8'b10010111;
DRAM[42844] = 8'b10011010;
DRAM[42845] = 8'b10011111;
DRAM[42846] = 8'b10100101;
DRAM[42847] = 8'b10101001;
DRAM[42848] = 8'b10101110;
DRAM[42849] = 8'b10110000;
DRAM[42850] = 8'b10110011;
DRAM[42851] = 8'b10110111;
DRAM[42852] = 8'b10111010;
DRAM[42853] = 8'b11000000;
DRAM[42854] = 8'b11000111;
DRAM[42855] = 8'b11001011;
DRAM[42856] = 8'b11000100;
DRAM[42857] = 8'b11001001;
DRAM[42858] = 8'b11001110;
DRAM[42859] = 8'b11001111;
DRAM[42860] = 8'b11001110;
DRAM[42861] = 8'b11001100;
DRAM[42862] = 8'b11001101;
DRAM[42863] = 8'b11001111;
DRAM[42864] = 8'b11010000;
DRAM[42865] = 8'b11001100;
DRAM[42866] = 8'b11001100;
DRAM[42867] = 8'b11000101;
DRAM[42868] = 8'b10110111;
DRAM[42869] = 8'b10110011;
DRAM[42870] = 8'b10101111;
DRAM[42871] = 8'b10100011;
DRAM[42872] = 8'b10100001;
DRAM[42873] = 8'b10011011;
DRAM[42874] = 8'b10010110;
DRAM[42875] = 8'b10010110;
DRAM[42876] = 8'b10011010;
DRAM[42877] = 8'b10011111;
DRAM[42878] = 8'b10100010;
DRAM[42879] = 8'b10100100;
DRAM[42880] = 8'b10011001;
DRAM[42881] = 8'b10001010;
DRAM[42882] = 8'b1110011;
DRAM[42883] = 8'b1100001;
DRAM[42884] = 8'b1011101;
DRAM[42885] = 8'b1011010;
DRAM[42886] = 8'b1000111;
DRAM[42887] = 8'b110000;
DRAM[42888] = 8'b11110;
DRAM[42889] = 8'b101;
DRAM[42890] = 8'b0;
DRAM[42891] = 8'b111;
DRAM[42892] = 8'b100;
DRAM[42893] = 8'b0;
DRAM[42894] = 8'b0;
DRAM[42895] = 8'b0;
DRAM[42896] = 8'b0;
DRAM[42897] = 8'b0;
DRAM[42898] = 8'b0;
DRAM[42899] = 8'b0;
DRAM[42900] = 8'b0;
DRAM[42901] = 8'b0;
DRAM[42902] = 8'b0;
DRAM[42903] = 8'b0;
DRAM[42904] = 8'b11;
DRAM[42905] = 8'b10;
DRAM[42906] = 8'b10;
DRAM[42907] = 8'b10;
DRAM[42908] = 8'b11;
DRAM[42909] = 8'b11;
DRAM[42910] = 8'b10;
DRAM[42911] = 8'b0;
DRAM[42912] = 8'b11100;
DRAM[42913] = 8'b110010;
DRAM[42914] = 8'b1001100;
DRAM[42915] = 8'b1010110;
DRAM[42916] = 8'b1011100;
DRAM[42917] = 8'b1110101;
DRAM[42918] = 8'b10001111;
DRAM[42919] = 8'b10010100;
DRAM[42920] = 8'b10010100;
DRAM[42921] = 8'b10011000;
DRAM[42922] = 8'b10100001;
DRAM[42923] = 8'b10101101;
DRAM[42924] = 8'b10110100;
DRAM[42925] = 8'b10111010;
DRAM[42926] = 8'b11000100;
DRAM[42927] = 8'b11001111;
DRAM[42928] = 8'b11011000;
DRAM[42929] = 8'b11101000;
DRAM[42930] = 8'b11101101;
DRAM[42931] = 8'b11011111;
DRAM[42932] = 8'b11010101;
DRAM[42933] = 8'b11010111;
DRAM[42934] = 8'b11010101;
DRAM[42935] = 8'b11001011;
DRAM[42936] = 8'b11011100;
DRAM[42937] = 8'b11011101;
DRAM[42938] = 8'b11100011;
DRAM[42939] = 8'b11010001;
DRAM[42940] = 8'b11001010;
DRAM[42941] = 8'b11010011;
DRAM[42942] = 8'b11001101;
DRAM[42943] = 8'b11010001;
DRAM[42944] = 8'b11010010;
DRAM[42945] = 8'b11010100;
DRAM[42946] = 8'b11010000;
DRAM[42947] = 8'b11000100;
DRAM[42948] = 8'b10110100;
DRAM[42949] = 8'b10101110;
DRAM[42950] = 8'b10110110;
DRAM[42951] = 8'b11000011;
DRAM[42952] = 8'b10110111;
DRAM[42953] = 8'b11000100;
DRAM[42954] = 8'b11001100;
DRAM[42955] = 8'b11000010;
DRAM[42956] = 8'b10101011;
DRAM[42957] = 8'b10011011;
DRAM[42958] = 8'b10011011;
DRAM[42959] = 8'b10100010;
DRAM[42960] = 8'b10011010;
DRAM[42961] = 8'b10011001;
DRAM[42962] = 8'b10011001;
DRAM[42963] = 8'b10011010;
DRAM[42964] = 8'b10011010;
DRAM[42965] = 8'b10011000;
DRAM[42966] = 8'b10010100;
DRAM[42967] = 8'b10010000;
DRAM[42968] = 8'b10010001;
DRAM[42969] = 8'b10010011;
DRAM[42970] = 8'b10010110;
DRAM[42971] = 8'b10011001;
DRAM[42972] = 8'b10011010;
DRAM[42973] = 8'b10011010;
DRAM[42974] = 8'b10011001;
DRAM[42975] = 8'b10011001;
DRAM[42976] = 8'b10000110;
DRAM[42977] = 8'b10000101;
DRAM[42978] = 8'b10000100;
DRAM[42979] = 8'b10000100;
DRAM[42980] = 8'b10000100;
DRAM[42981] = 8'b10000011;
DRAM[42982] = 8'b10000000;
DRAM[42983] = 8'b1111110;
DRAM[42984] = 8'b1111100;
DRAM[42985] = 8'b1111100;
DRAM[42986] = 8'b1111011;
DRAM[42987] = 8'b1111011;
DRAM[42988] = 8'b1111011;
DRAM[42989] = 8'b1111100;
DRAM[42990] = 8'b1111101;
DRAM[42991] = 8'b1111101;
DRAM[42992] = 8'b10000000;
DRAM[42993] = 8'b10000000;
DRAM[42994] = 8'b10000000;
DRAM[42995] = 8'b10000001;
DRAM[42996] = 8'b10000010;
DRAM[42997] = 8'b10000011;
DRAM[42998] = 8'b10000101;
DRAM[42999] = 8'b10000110;
DRAM[43000] = 8'b10000011;
DRAM[43001] = 8'b10000010;
DRAM[43002] = 8'b10000011;
DRAM[43003] = 8'b10000110;
DRAM[43004] = 8'b10001000;
DRAM[43005] = 8'b10001000;
DRAM[43006] = 8'b10000110;
DRAM[43007] = 8'b10000100;
DRAM[43008] = 8'b10010101;
DRAM[43009] = 8'b10010101;
DRAM[43010] = 8'b10010110;
DRAM[43011] = 8'b10010110;
DRAM[43012] = 8'b10010110;
DRAM[43013] = 8'b10010111;
DRAM[43014] = 8'b10010111;
DRAM[43015] = 8'b10010111;
DRAM[43016] = 8'b10011001;
DRAM[43017] = 8'b10011010;
DRAM[43018] = 8'b10011011;
DRAM[43019] = 8'b10011101;
DRAM[43020] = 8'b10011101;
DRAM[43021] = 8'b10011110;
DRAM[43022] = 8'b10011110;
DRAM[43023] = 8'b10011101;
DRAM[43024] = 8'b10011111;
DRAM[43025] = 8'b10100000;
DRAM[43026] = 8'b10100000;
DRAM[43027] = 8'b10100000;
DRAM[43028] = 8'b10100000;
DRAM[43029] = 8'b10100000;
DRAM[43030] = 8'b10100001;
DRAM[43031] = 8'b10100001;
DRAM[43032] = 8'b10100010;
DRAM[43033] = 8'b10100010;
DRAM[43034] = 8'b10100010;
DRAM[43035] = 8'b10100010;
DRAM[43036] = 8'b10100011;
DRAM[43037] = 8'b10100100;
DRAM[43038] = 8'b10100101;
DRAM[43039] = 8'b10100110;
DRAM[43040] = 8'b10100010;
DRAM[43041] = 8'b10100101;
DRAM[43042] = 8'b10100110;
DRAM[43043] = 8'b10100011;
DRAM[43044] = 8'b10100111;
DRAM[43045] = 8'b10111011;
DRAM[43046] = 8'b11011100;
DRAM[43047] = 8'b11110110;
DRAM[43048] = 8'b11111101;
DRAM[43049] = 8'b11111101;
DRAM[43050] = 8'b11111101;
DRAM[43051] = 8'b11111110;
DRAM[43052] = 8'b11111110;
DRAM[43053] = 8'b11111111;
DRAM[43054] = 8'b11111111;
DRAM[43055] = 8'b11111111;
DRAM[43056] = 8'b11111101;
DRAM[43057] = 8'b11111101;
DRAM[43058] = 8'b11111101;
DRAM[43059] = 8'b11111110;
DRAM[43060] = 8'b11111110;
DRAM[43061] = 8'b11111111;
DRAM[43062] = 8'b11111111;
DRAM[43063] = 8'b11111111;
DRAM[43064] = 8'b11111111;
DRAM[43065] = 8'b11111011;
DRAM[43066] = 8'b11110111;
DRAM[43067] = 8'b11110111;
DRAM[43068] = 8'b11110111;
DRAM[43069] = 8'b11110101;
DRAM[43070] = 8'b11110000;
DRAM[43071] = 8'b11101011;
DRAM[43072] = 8'b11101011;
DRAM[43073] = 8'b11100100;
DRAM[43074] = 8'b11011010;
DRAM[43075] = 8'b11010010;
DRAM[43076] = 8'b11001101;
DRAM[43077] = 8'b11001011;
DRAM[43078] = 8'b11001010;
DRAM[43079] = 8'b11001001;
DRAM[43080] = 8'b11001001;
DRAM[43081] = 8'b10111110;
DRAM[43082] = 8'b10110111;
DRAM[43083] = 8'b10111000;
DRAM[43084] = 8'b10110110;
DRAM[43085] = 8'b10101110;
DRAM[43086] = 8'b10100111;
DRAM[43087] = 8'b10100101;
DRAM[43088] = 8'b10011110;
DRAM[43089] = 8'b10011010;
DRAM[43090] = 8'b10010110;
DRAM[43091] = 8'b10011000;
DRAM[43092] = 8'b10011011;
DRAM[43093] = 8'b10011011;
DRAM[43094] = 8'b10010101;
DRAM[43095] = 8'b10001111;
DRAM[43096] = 8'b10001011;
DRAM[43097] = 8'b10010100;
DRAM[43098] = 8'b10011101;
DRAM[43099] = 8'b10011110;
DRAM[43100] = 8'b10011100;
DRAM[43101] = 8'b10011111;
DRAM[43102] = 8'b10101001;
DRAM[43103] = 8'b10110011;
DRAM[43104] = 8'b10101011;
DRAM[43105] = 8'b10101001;
DRAM[43106] = 8'b10101010;
DRAM[43107] = 8'b10101111;
DRAM[43108] = 8'b10110000;
DRAM[43109] = 8'b10110000;
DRAM[43110] = 8'b10110111;
DRAM[43111] = 8'b11000001;
DRAM[43112] = 8'b10110110;
DRAM[43113] = 8'b10111110;
DRAM[43114] = 8'b11000000;
DRAM[43115] = 8'b10111100;
DRAM[43116] = 8'b11000000;
DRAM[43117] = 8'b11001011;
DRAM[43118] = 8'b11001110;
DRAM[43119] = 8'b11001000;
DRAM[43120] = 8'b11001010;
DRAM[43121] = 8'b11001101;
DRAM[43122] = 8'b11001111;
DRAM[43123] = 8'b11001111;
DRAM[43124] = 8'b11001111;
DRAM[43125] = 8'b11001010;
DRAM[43126] = 8'b10111100;
DRAM[43127] = 8'b10101111;
DRAM[43128] = 8'b10101011;
DRAM[43129] = 8'b10011100;
DRAM[43130] = 8'b10001111;
DRAM[43131] = 8'b10010001;
DRAM[43132] = 8'b10011011;
DRAM[43133] = 8'b10100100;
DRAM[43134] = 8'b10101001;
DRAM[43135] = 8'b10101101;
DRAM[43136] = 8'b10011010;
DRAM[43137] = 8'b10001111;
DRAM[43138] = 8'b1111010;
DRAM[43139] = 8'b1101000;
DRAM[43140] = 8'b1100101;
DRAM[43141] = 8'b1100001;
DRAM[43142] = 8'b1001000;
DRAM[43143] = 8'b101001;
DRAM[43144] = 8'b11001;
DRAM[43145] = 8'b1101;
DRAM[43146] = 8'b10;
DRAM[43147] = 8'b0;
DRAM[43148] = 8'b0;
DRAM[43149] = 8'b0;
DRAM[43150] = 8'b0;
DRAM[43151] = 8'b10;
DRAM[43152] = 8'b0;
DRAM[43153] = 8'b0;
DRAM[43154] = 8'b0;
DRAM[43155] = 8'b0;
DRAM[43156] = 8'b0;
DRAM[43157] = 8'b0;
DRAM[43158] = 8'b0;
DRAM[43159] = 8'b0;
DRAM[43160] = 8'b0;
DRAM[43161] = 8'b0;
DRAM[43162] = 8'b0;
DRAM[43163] = 8'b0;
DRAM[43164] = 8'b0;
DRAM[43165] = 8'b0;
DRAM[43166] = 8'b0;
DRAM[43167] = 8'b1;
DRAM[43168] = 8'b1101;
DRAM[43169] = 8'b101100;
DRAM[43170] = 8'b1000111;
DRAM[43171] = 8'b1011001;
DRAM[43172] = 8'b1101000;
DRAM[43173] = 8'b1101110;
DRAM[43174] = 8'b1111001;
DRAM[43175] = 8'b10001011;
DRAM[43176] = 8'b10001100;
DRAM[43177] = 8'b10100000;
DRAM[43178] = 8'b10101011;
DRAM[43179] = 8'b10100110;
DRAM[43180] = 8'b10101010;
DRAM[43181] = 8'b10111101;
DRAM[43182] = 8'b11001011;
DRAM[43183] = 8'b11001011;
DRAM[43184] = 8'b11001101;
DRAM[43185] = 8'b11101001;
DRAM[43186] = 8'b11100110;
DRAM[43187] = 8'b11010100;
DRAM[43188] = 8'b11010100;
DRAM[43189] = 8'b11010001;
DRAM[43190] = 8'b11001001;
DRAM[43191] = 8'b11001110;
DRAM[43192] = 8'b11101111;
DRAM[43193] = 8'b11011011;
DRAM[43194] = 8'b10100101;
DRAM[43195] = 8'b10110011;
DRAM[43196] = 8'b11010011;
DRAM[43197] = 8'b11010000;
DRAM[43198] = 8'b11011111;
DRAM[43199] = 8'b11100111;
DRAM[43200] = 8'b11100000;
DRAM[43201] = 8'b11000100;
DRAM[43202] = 8'b10110000;
DRAM[43203] = 8'b10111001;
DRAM[43204] = 8'b11001011;
DRAM[43205] = 8'b11001111;
DRAM[43206] = 8'b11000000;
DRAM[43207] = 8'b10110001;
DRAM[43208] = 8'b10110101;
DRAM[43209] = 8'b10101111;
DRAM[43210] = 8'b10110100;
DRAM[43211] = 8'b11000100;
DRAM[43212] = 8'b11001000;
DRAM[43213] = 8'b10110110;
DRAM[43214] = 8'b10011111;
DRAM[43215] = 8'b10010010;
DRAM[43216] = 8'b10100001;
DRAM[43217] = 8'b10011011;
DRAM[43218] = 8'b10011001;
DRAM[43219] = 8'b10011100;
DRAM[43220] = 8'b10011100;
DRAM[43221] = 8'b10010110;
DRAM[43222] = 8'b10010000;
DRAM[43223] = 8'b10001110;
DRAM[43224] = 8'b10010010;
DRAM[43225] = 8'b10010000;
DRAM[43226] = 8'b10001111;
DRAM[43227] = 8'b10001111;
DRAM[43228] = 8'b10001111;
DRAM[43229] = 8'b10001110;
DRAM[43230] = 8'b10001011;
DRAM[43231] = 8'b10001001;
DRAM[43232] = 8'b10000111;
DRAM[43233] = 8'b10000101;
DRAM[43234] = 8'b10000011;
DRAM[43235] = 8'b10000010;
DRAM[43236] = 8'b10000010;
DRAM[43237] = 8'b10000001;
DRAM[43238] = 8'b1111111;
DRAM[43239] = 8'b1111101;
DRAM[43240] = 8'b1111011;
DRAM[43241] = 8'b1111100;
DRAM[43242] = 8'b1111101;
DRAM[43243] = 8'b1111101;
DRAM[43244] = 8'b1111110;
DRAM[43245] = 8'b1111110;
DRAM[43246] = 8'b1111110;
DRAM[43247] = 8'b1111101;
DRAM[43248] = 8'b10000000;
DRAM[43249] = 8'b10000001;
DRAM[43250] = 8'b10000010;
DRAM[43251] = 8'b10000100;
DRAM[43252] = 8'b10000101;
DRAM[43253] = 8'b10000110;
DRAM[43254] = 8'b10000111;
DRAM[43255] = 8'b10000111;
DRAM[43256] = 8'b10000101;
DRAM[43257] = 8'b10000101;
DRAM[43258] = 8'b10000101;
DRAM[43259] = 8'b10000101;
DRAM[43260] = 8'b10000101;
DRAM[43261] = 8'b10000101;
DRAM[43262] = 8'b10000101;
DRAM[43263] = 8'b10000101;
DRAM[43264] = 8'b10010101;
DRAM[43265] = 8'b10010101;
DRAM[43266] = 8'b10010101;
DRAM[43267] = 8'b10010110;
DRAM[43268] = 8'b10010110;
DRAM[43269] = 8'b10010110;
DRAM[43270] = 8'b10010111;
DRAM[43271] = 8'b10010111;
DRAM[43272] = 8'b10011000;
DRAM[43273] = 8'b10011001;
DRAM[43274] = 8'b10011010;
DRAM[43275] = 8'b10011100;
DRAM[43276] = 8'b10011100;
DRAM[43277] = 8'b10011101;
DRAM[43278] = 8'b10011101;
DRAM[43279] = 8'b10011101;
DRAM[43280] = 8'b10011111;
DRAM[43281] = 8'b10011111;
DRAM[43282] = 8'b10011111;
DRAM[43283] = 8'b10100000;
DRAM[43284] = 8'b10100000;
DRAM[43285] = 8'b10100000;
DRAM[43286] = 8'b10100000;
DRAM[43287] = 8'b10100001;
DRAM[43288] = 8'b10100010;
DRAM[43289] = 8'b10100001;
DRAM[43290] = 8'b10100001;
DRAM[43291] = 8'b10100010;
DRAM[43292] = 8'b10100010;
DRAM[43293] = 8'b10100100;
DRAM[43294] = 8'b10100101;
DRAM[43295] = 8'b10100110;
DRAM[43296] = 8'b10100011;
DRAM[43297] = 8'b10100110;
DRAM[43298] = 8'b10101001;
DRAM[43299] = 8'b10101100;
DRAM[43300] = 8'b10110110;
DRAM[43301] = 8'b11001010;
DRAM[43302] = 8'b11100100;
DRAM[43303] = 8'b11110111;
DRAM[43304] = 8'b11111101;
DRAM[43305] = 8'b11111101;
DRAM[43306] = 8'b11111101;
DRAM[43307] = 8'b11111110;
DRAM[43308] = 8'b11111110;
DRAM[43309] = 8'b11111111;
DRAM[43310] = 8'b11111111;
DRAM[43311] = 8'b11111111;
DRAM[43312] = 8'b11111101;
DRAM[43313] = 8'b11111101;
DRAM[43314] = 8'b11111101;
DRAM[43315] = 8'b11111110;
DRAM[43316] = 8'b11111110;
DRAM[43317] = 8'b11111111;
DRAM[43318] = 8'b11111111;
DRAM[43319] = 8'b11111111;
DRAM[43320] = 8'b11111100;
DRAM[43321] = 8'b11111100;
DRAM[43322] = 8'b11111011;
DRAM[43323] = 8'b11111000;
DRAM[43324] = 8'b11110101;
DRAM[43325] = 8'b11110001;
DRAM[43326] = 8'b11101111;
DRAM[43327] = 8'b11101110;
DRAM[43328] = 8'b11100010;
DRAM[43329] = 8'b11100000;
DRAM[43330] = 8'b11011110;
DRAM[43331] = 8'b11011011;
DRAM[43332] = 8'b11010110;
DRAM[43333] = 8'b11001101;
DRAM[43334] = 8'b11000011;
DRAM[43335] = 8'b10111100;
DRAM[43336] = 8'b11001101;
DRAM[43337] = 8'b11000100;
DRAM[43338] = 8'b10111101;
DRAM[43339] = 8'b10111011;
DRAM[43340] = 8'b10110110;
DRAM[43341] = 8'b10101100;
DRAM[43342] = 8'b10100100;
DRAM[43343] = 8'b10100010;
DRAM[43344] = 8'b10100111;
DRAM[43345] = 8'b10100110;
DRAM[43346] = 8'b10100100;
DRAM[43347] = 8'b10100000;
DRAM[43348] = 8'b10011010;
DRAM[43349] = 8'b10010001;
DRAM[43350] = 8'b10001000;
DRAM[43351] = 8'b10000011;
DRAM[43352] = 8'b10001110;
DRAM[43353] = 8'b10010000;
DRAM[43354] = 8'b10010010;
DRAM[43355] = 8'b10010001;
DRAM[43356] = 8'b10010000;
DRAM[43357] = 8'b10010001;
DRAM[43358] = 8'b10010110;
DRAM[43359] = 8'b10011010;
DRAM[43360] = 8'b10110000;
DRAM[43361] = 8'b10101110;
DRAM[43362] = 8'b10110001;
DRAM[43363] = 8'b10110110;
DRAM[43364] = 8'b10110110;
DRAM[43365] = 8'b10110100;
DRAM[43366] = 8'b10111000;
DRAM[43367] = 8'b11000000;
DRAM[43368] = 8'b10110111;
DRAM[43369] = 8'b10111011;
DRAM[43370] = 8'b10111001;
DRAM[43371] = 8'b10110110;
DRAM[43372] = 8'b10111101;
DRAM[43373] = 8'b11001010;
DRAM[43374] = 8'b11001100;
DRAM[43375] = 8'b11000101;
DRAM[43376] = 8'b11001000;
DRAM[43377] = 8'b11001101;
DRAM[43378] = 8'b11010010;
DRAM[43379] = 8'b11010100;
DRAM[43380] = 8'b11010100;
DRAM[43381] = 8'b11001100;
DRAM[43382] = 8'b10111011;
DRAM[43383] = 8'b10101011;
DRAM[43384] = 8'b10110100;
DRAM[43385] = 8'b10100110;
DRAM[43386] = 8'b10011010;
DRAM[43387] = 8'b10011011;
DRAM[43388] = 8'b10100000;
DRAM[43389] = 8'b10100011;
DRAM[43390] = 8'b10100100;
DRAM[43391] = 8'b10100100;
DRAM[43392] = 8'b10010101;
DRAM[43393] = 8'b10000010;
DRAM[43394] = 8'b1110101;
DRAM[43395] = 8'b1110110;
DRAM[43396] = 8'b1101111;
DRAM[43397] = 8'b1011001;
DRAM[43398] = 8'b1000100;
DRAM[43399] = 8'b111100;
DRAM[43400] = 8'b100010;
DRAM[43401] = 8'b10010;
DRAM[43402] = 8'b10;
DRAM[43403] = 8'b0;
DRAM[43404] = 8'b11;
DRAM[43405] = 8'b11;
DRAM[43406] = 8'b1;
DRAM[43407] = 8'b0;
DRAM[43408] = 8'b0;
DRAM[43409] = 8'b0;
DRAM[43410] = 8'b0;
DRAM[43411] = 8'b0;
DRAM[43412] = 8'b0;
DRAM[43413] = 8'b0;
DRAM[43414] = 8'b0;
DRAM[43415] = 8'b0;
DRAM[43416] = 8'b0;
DRAM[43417] = 8'b0;
DRAM[43418] = 8'b0;
DRAM[43419] = 8'b0;
DRAM[43420] = 8'b0;
DRAM[43421] = 8'b10;
DRAM[43422] = 8'b100;
DRAM[43423] = 8'b101;
DRAM[43424] = 8'b11000;
DRAM[43425] = 8'b110010;
DRAM[43426] = 8'b1000111;
DRAM[43427] = 8'b1010101;
DRAM[43428] = 8'b1100010;
DRAM[43429] = 8'b1101000;
DRAM[43430] = 8'b1110010;
DRAM[43431] = 8'b10000011;
DRAM[43432] = 8'b10010100;
DRAM[43433] = 8'b10100011;
DRAM[43434] = 8'b10101110;
DRAM[43435] = 8'b10110001;
DRAM[43436] = 8'b10110110;
DRAM[43437] = 8'b10111111;
DRAM[43438] = 8'b11000001;
DRAM[43439] = 8'b10111101;
DRAM[43440] = 8'b11010001;
DRAM[43441] = 8'b11100110;
DRAM[43442] = 8'b11100111;
DRAM[43443] = 8'b11011101;
DRAM[43444] = 8'b11011010;
DRAM[43445] = 8'b11001110;
DRAM[43446] = 8'b11001011;
DRAM[43447] = 8'b11011011;
DRAM[43448] = 8'b11010111;
DRAM[43449] = 8'b11011000;
DRAM[43450] = 8'b10111000;
DRAM[43451] = 8'b10101000;
DRAM[43452] = 8'b10110110;
DRAM[43453] = 8'b11001110;
DRAM[43454] = 8'b11100010;
DRAM[43455] = 8'b11011111;
DRAM[43456] = 8'b11101011;
DRAM[43457] = 8'b11101001;
DRAM[43458] = 8'b11100010;
DRAM[43459] = 8'b11010000;
DRAM[43460] = 8'b10110111;
DRAM[43461] = 8'b10101000;
DRAM[43462] = 8'b10110000;
DRAM[43463] = 8'b11000001;
DRAM[43464] = 8'b10110100;
DRAM[43465] = 8'b10101101;
DRAM[43466] = 8'b10011111;
DRAM[43467] = 8'b10011010;
DRAM[43468] = 8'b10101100;
DRAM[43469] = 8'b11000000;
DRAM[43470] = 8'b10111100;
DRAM[43471] = 8'b10101001;
DRAM[43472] = 8'b10100000;
DRAM[43473] = 8'b10011010;
DRAM[43474] = 8'b10010111;
DRAM[43475] = 8'b10011001;
DRAM[43476] = 8'b10011001;
DRAM[43477] = 8'b10010110;
DRAM[43478] = 8'b10010011;
DRAM[43479] = 8'b10010100;
DRAM[43480] = 8'b10010001;
DRAM[43481] = 8'b10010000;
DRAM[43482] = 8'b10001110;
DRAM[43483] = 8'b10001110;
DRAM[43484] = 8'b10001111;
DRAM[43485] = 8'b10001110;
DRAM[43486] = 8'b10001011;
DRAM[43487] = 8'b10001001;
DRAM[43488] = 8'b10000111;
DRAM[43489] = 8'b10000100;
DRAM[43490] = 8'b10000010;
DRAM[43491] = 8'b10000001;
DRAM[43492] = 8'b10000001;
DRAM[43493] = 8'b1111111;
DRAM[43494] = 8'b1111101;
DRAM[43495] = 8'b1111011;
DRAM[43496] = 8'b1111001;
DRAM[43497] = 8'b1111010;
DRAM[43498] = 8'b1111011;
DRAM[43499] = 8'b1111101;
DRAM[43500] = 8'b1111110;
DRAM[43501] = 8'b1111111;
DRAM[43502] = 8'b10000000;
DRAM[43503] = 8'b10000000;
DRAM[43504] = 8'b10000000;
DRAM[43505] = 8'b10000001;
DRAM[43506] = 8'b10000011;
DRAM[43507] = 8'b10000100;
DRAM[43508] = 8'b10000110;
DRAM[43509] = 8'b10000110;
DRAM[43510] = 8'b10000111;
DRAM[43511] = 8'b10000111;
DRAM[43512] = 8'b10000101;
DRAM[43513] = 8'b10000101;
DRAM[43514] = 8'b10000101;
DRAM[43515] = 8'b10000101;
DRAM[43516] = 8'b10000101;
DRAM[43517] = 8'b10000101;
DRAM[43518] = 8'b10000101;
DRAM[43519] = 8'b10000101;
DRAM[43520] = 8'b10010100;
DRAM[43521] = 8'b10010100;
DRAM[43522] = 8'b10010101;
DRAM[43523] = 8'b10010101;
DRAM[43524] = 8'b10010101;
DRAM[43525] = 8'b10010110;
DRAM[43526] = 8'b10010110;
DRAM[43527] = 8'b10010110;
DRAM[43528] = 8'b10010111;
DRAM[43529] = 8'b10011000;
DRAM[43530] = 8'b10011001;
DRAM[43531] = 8'b10011010;
DRAM[43532] = 8'b10011011;
DRAM[43533] = 8'b10011011;
DRAM[43534] = 8'b10011011;
DRAM[43535] = 8'b10011011;
DRAM[43536] = 8'b10011110;
DRAM[43537] = 8'b10011110;
DRAM[43538] = 8'b10011110;
DRAM[43539] = 8'b10011111;
DRAM[43540] = 8'b10011111;
DRAM[43541] = 8'b10100000;
DRAM[43542] = 8'b10100000;
DRAM[43543] = 8'b10100000;
DRAM[43544] = 8'b10100001;
DRAM[43545] = 8'b10100001;
DRAM[43546] = 8'b10100001;
DRAM[43547] = 8'b10100001;
DRAM[43548] = 8'b10100010;
DRAM[43549] = 8'b10100011;
DRAM[43550] = 8'b10100101;
DRAM[43551] = 8'b10100101;
DRAM[43552] = 8'b10100101;
DRAM[43553] = 8'b10100111;
DRAM[43554] = 8'b10101011;
DRAM[43555] = 8'b10110101;
DRAM[43556] = 8'b11000101;
DRAM[43557] = 8'b11011010;
DRAM[43558] = 8'b11101101;
DRAM[43559] = 8'b11111010;
DRAM[43560] = 8'b11111101;
DRAM[43561] = 8'b11111101;
DRAM[43562] = 8'b11111101;
DRAM[43563] = 8'b11111110;
DRAM[43564] = 8'b11111110;
DRAM[43565] = 8'b11111111;
DRAM[43566] = 8'b11111111;
DRAM[43567] = 8'b11111111;
DRAM[43568] = 8'b11111101;
DRAM[43569] = 8'b11111101;
DRAM[43570] = 8'b11111110;
DRAM[43571] = 8'b11111110;
DRAM[43572] = 8'b11111110;
DRAM[43573] = 8'b11111110;
DRAM[43574] = 8'b11111111;
DRAM[43575] = 8'b11111111;
DRAM[43576] = 8'b11111001;
DRAM[43577] = 8'b11111100;
DRAM[43578] = 8'b11111101;
DRAM[43579] = 8'b11111001;
DRAM[43580] = 8'b11110011;
DRAM[43581] = 8'b11101110;
DRAM[43582] = 8'b11101110;
DRAM[43583] = 8'b11110000;
DRAM[43584] = 8'b11100110;
DRAM[43585] = 8'b11100001;
DRAM[43586] = 8'b11011010;
DRAM[43587] = 8'b11010100;
DRAM[43588] = 8'b11001111;
DRAM[43589] = 8'b11001011;
DRAM[43590] = 8'b11001000;
DRAM[43591] = 8'b11000101;
DRAM[43592] = 8'b11000101;
DRAM[43593] = 8'b11000001;
DRAM[43594] = 8'b11000000;
DRAM[43595] = 8'b10111111;
DRAM[43596] = 8'b10111011;
DRAM[43597] = 8'b10110100;
DRAM[43598] = 8'b10101111;
DRAM[43599] = 8'b10101111;
DRAM[43600] = 8'b10101000;
DRAM[43601] = 8'b10101001;
DRAM[43602] = 8'b10100111;
DRAM[43603] = 8'b10100001;
DRAM[43604] = 8'b10011000;
DRAM[43605] = 8'b10010001;
DRAM[43606] = 8'b10001110;
DRAM[43607] = 8'b10001101;
DRAM[43608] = 8'b10010000;
DRAM[43609] = 8'b10001101;
DRAM[43610] = 8'b10001010;
DRAM[43611] = 8'b10001010;
DRAM[43612] = 8'b10001100;
DRAM[43613] = 8'b10001111;
DRAM[43614] = 8'b10010001;
DRAM[43615] = 8'b10010010;
DRAM[43616] = 8'b10100000;
DRAM[43617] = 8'b10100010;
DRAM[43618] = 8'b10100111;
DRAM[43619] = 8'b10101110;
DRAM[43620] = 8'b10101111;
DRAM[43621] = 8'b10101101;
DRAM[43622] = 8'b10101101;
DRAM[43623] = 8'b10110001;
DRAM[43624] = 8'b10101111;
DRAM[43625] = 8'b10101111;
DRAM[43626] = 8'b10101100;
DRAM[43627] = 8'b10101011;
DRAM[43628] = 8'b10110110;
DRAM[43629] = 8'b11000101;
DRAM[43630] = 8'b11000111;
DRAM[43631] = 8'b11000000;
DRAM[43632] = 8'b11001111;
DRAM[43633] = 8'b11010011;
DRAM[43634] = 8'b11010101;
DRAM[43635] = 8'b11010010;
DRAM[43636] = 8'b11001100;
DRAM[43637] = 8'b11000010;
DRAM[43638] = 8'b10110100;
DRAM[43639] = 8'b10100111;
DRAM[43640] = 8'b10110111;
DRAM[43641] = 8'b10101011;
DRAM[43642] = 8'b10100010;
DRAM[43643] = 8'b10100011;
DRAM[43644] = 8'b10100101;
DRAM[43645] = 8'b10100010;
DRAM[43646] = 8'b10011101;
DRAM[43647] = 8'b10011010;
DRAM[43648] = 8'b10000110;
DRAM[43649] = 8'b1111000;
DRAM[43650] = 8'b1101111;
DRAM[43651] = 8'b1101101;
DRAM[43652] = 8'b1100001;
DRAM[43653] = 8'b1001101;
DRAM[43654] = 8'b1000011;
DRAM[43655] = 8'b1000101;
DRAM[43656] = 8'b101101;
DRAM[43657] = 8'b11001;
DRAM[43658] = 8'b110;
DRAM[43659] = 8'b10;
DRAM[43660] = 8'b110;
DRAM[43661] = 8'b110;
DRAM[43662] = 8'b10;
DRAM[43663] = 8'b0;
DRAM[43664] = 8'b0;
DRAM[43665] = 8'b0;
DRAM[43666] = 8'b0;
DRAM[43667] = 8'b0;
DRAM[43668] = 8'b0;
DRAM[43669] = 8'b0;
DRAM[43670] = 8'b0;
DRAM[43671] = 8'b0;
DRAM[43672] = 8'b0;
DRAM[43673] = 8'b0;
DRAM[43674] = 8'b0;
DRAM[43675] = 8'b0;
DRAM[43676] = 8'b1;
DRAM[43677] = 8'b101;
DRAM[43678] = 8'b1001;
DRAM[43679] = 8'b1100;
DRAM[43680] = 8'b101000;
DRAM[43681] = 8'b111011;
DRAM[43682] = 8'b1001001;
DRAM[43683] = 8'b1010101;
DRAM[43684] = 8'b1100100;
DRAM[43685] = 8'b1101011;
DRAM[43686] = 8'b1110100;
DRAM[43687] = 8'b10000011;
DRAM[43688] = 8'b10011011;
DRAM[43689] = 8'b10100001;
DRAM[43690] = 8'b10101010;
DRAM[43691] = 8'b10110100;
DRAM[43692] = 8'b10111011;
DRAM[43693] = 8'b10111110;
DRAM[43694] = 8'b10111101;
DRAM[43695] = 8'b10111011;
DRAM[43696] = 8'b11010100;
DRAM[43697] = 8'b11100000;
DRAM[43698] = 8'b11100101;
DRAM[43699] = 8'b11100100;
DRAM[43700] = 8'b11011111;
DRAM[43701] = 8'b11010001;
DRAM[43702] = 8'b11010011;
DRAM[43703] = 8'b11101001;
DRAM[43704] = 8'b11000111;
DRAM[43705] = 8'b10101110;
DRAM[43706] = 8'b10101110;
DRAM[43707] = 8'b10110010;
DRAM[43708] = 8'b10111100;
DRAM[43709] = 8'b11001111;
DRAM[43710] = 8'b11011010;
DRAM[43711] = 8'b11100111;
DRAM[43712] = 8'b11100100;
DRAM[43713] = 8'b11010111;
DRAM[43714] = 8'b11010001;
DRAM[43715] = 8'b11011000;
DRAM[43716] = 8'b11011111;
DRAM[43717] = 8'b11010011;
DRAM[43718] = 8'b10110111;
DRAM[43719] = 8'b10100001;
DRAM[43720] = 8'b10100100;
DRAM[43721] = 8'b10101011;
DRAM[43722] = 8'b10101001;
DRAM[43723] = 8'b10011110;
DRAM[43724] = 8'b10011110;
DRAM[43725] = 8'b10101011;
DRAM[43726] = 8'b10110011;
DRAM[43727] = 8'b10110001;
DRAM[43728] = 8'b10100011;
DRAM[43729] = 8'b10011100;
DRAM[43730] = 8'b10010111;
DRAM[43731] = 8'b10010111;
DRAM[43732] = 8'b10010110;
DRAM[43733] = 8'b10010011;
DRAM[43734] = 8'b10010010;
DRAM[43735] = 8'b10010100;
DRAM[43736] = 8'b10010000;
DRAM[43737] = 8'b10001111;
DRAM[43738] = 8'b10001110;
DRAM[43739] = 8'b10001101;
DRAM[43740] = 8'b10001110;
DRAM[43741] = 8'b10001101;
DRAM[43742] = 8'b10001010;
DRAM[43743] = 8'b10001000;
DRAM[43744] = 8'b10000110;
DRAM[43745] = 8'b10000100;
DRAM[43746] = 8'b10000001;
DRAM[43747] = 8'b10000000;
DRAM[43748] = 8'b1111111;
DRAM[43749] = 8'b1111110;
DRAM[43750] = 8'b1111011;
DRAM[43751] = 8'b1111001;
DRAM[43752] = 8'b1111000;
DRAM[43753] = 8'b1111001;
DRAM[43754] = 8'b1111010;
DRAM[43755] = 8'b1111100;
DRAM[43756] = 8'b1111111;
DRAM[43757] = 8'b10000000;
DRAM[43758] = 8'b10000010;
DRAM[43759] = 8'b10000011;
DRAM[43760] = 8'b10000001;
DRAM[43761] = 8'b10000010;
DRAM[43762] = 8'b10000011;
DRAM[43763] = 8'b10000101;
DRAM[43764] = 8'b10000110;
DRAM[43765] = 8'b10000110;
DRAM[43766] = 8'b10000111;
DRAM[43767] = 8'b10000110;
DRAM[43768] = 8'b10000110;
DRAM[43769] = 8'b10000110;
DRAM[43770] = 8'b10000110;
DRAM[43771] = 8'b10000110;
DRAM[43772] = 8'b10000110;
DRAM[43773] = 8'b10000110;
DRAM[43774] = 8'b10000110;
DRAM[43775] = 8'b10000110;
DRAM[43776] = 8'b10010011;
DRAM[43777] = 8'b10010100;
DRAM[43778] = 8'b10010100;
DRAM[43779] = 8'b10010100;
DRAM[43780] = 8'b10010101;
DRAM[43781] = 8'b10010101;
DRAM[43782] = 8'b10010101;
DRAM[43783] = 8'b10010101;
DRAM[43784] = 8'b10010101;
DRAM[43785] = 8'b10010110;
DRAM[43786] = 8'b10010111;
DRAM[43787] = 8'b10011001;
DRAM[43788] = 8'b10011010;
DRAM[43789] = 8'b10011010;
DRAM[43790] = 8'b10011010;
DRAM[43791] = 8'b10011010;
DRAM[43792] = 8'b10011101;
DRAM[43793] = 8'b10011101;
DRAM[43794] = 8'b10011101;
DRAM[43795] = 8'b10011110;
DRAM[43796] = 8'b10011111;
DRAM[43797] = 8'b10011111;
DRAM[43798] = 8'b10100000;
DRAM[43799] = 8'b10100000;
DRAM[43800] = 8'b10100001;
DRAM[43801] = 8'b10100001;
DRAM[43802] = 8'b10100001;
DRAM[43803] = 8'b10100001;
DRAM[43804] = 8'b10100010;
DRAM[43805] = 8'b10100011;
DRAM[43806] = 8'b10100100;
DRAM[43807] = 8'b10100101;
DRAM[43808] = 8'b10100111;
DRAM[43809] = 8'b10101000;
DRAM[43810] = 8'b10101101;
DRAM[43811] = 8'b10110111;
DRAM[43812] = 8'b11000111;
DRAM[43813] = 8'b11011101;
DRAM[43814] = 8'b11110001;
DRAM[43815] = 8'b11111101;
DRAM[43816] = 8'b11111101;
DRAM[43817] = 8'b11111101;
DRAM[43818] = 8'b11111101;
DRAM[43819] = 8'b11111110;
DRAM[43820] = 8'b11111110;
DRAM[43821] = 8'b11111111;
DRAM[43822] = 8'b11111111;
DRAM[43823] = 8'b11111111;
DRAM[43824] = 8'b11111110;
DRAM[43825] = 8'b11111110;
DRAM[43826] = 8'b11111110;
DRAM[43827] = 8'b11111110;
DRAM[43828] = 8'b11111110;
DRAM[43829] = 8'b11111110;
DRAM[43830] = 8'b11111110;
DRAM[43831] = 8'b11111110;
DRAM[43832] = 8'b11111001;
DRAM[43833] = 8'b11111011;
DRAM[43834] = 8'b11111011;
DRAM[43835] = 8'b11111000;
DRAM[43836] = 8'b11110011;
DRAM[43837] = 8'b11101111;
DRAM[43838] = 8'b11101101;
DRAM[43839] = 8'b11101110;
DRAM[43840] = 8'b11100110;
DRAM[43841] = 8'b11100000;
DRAM[43842] = 8'b11011000;
DRAM[43843] = 8'b11010001;
DRAM[43844] = 8'b11001111;
DRAM[43845] = 8'b11010000;
DRAM[43846] = 8'b11010000;
DRAM[43847] = 8'b11010001;
DRAM[43848] = 8'b10111011;
DRAM[43849] = 8'b10111100;
DRAM[43850] = 8'b10111110;
DRAM[43851] = 8'b10111110;
DRAM[43852] = 8'b10111010;
DRAM[43853] = 8'b10110110;
DRAM[43854] = 8'b10110100;
DRAM[43855] = 8'b10110100;
DRAM[43856] = 8'b10101011;
DRAM[43857] = 8'b10101000;
DRAM[43858] = 8'b10100001;
DRAM[43859] = 8'b10011011;
DRAM[43860] = 8'b10010110;
DRAM[43861] = 8'b10010110;
DRAM[43862] = 8'b10011001;
DRAM[43863] = 8'b10011011;
DRAM[43864] = 8'b10001010;
DRAM[43865] = 8'b10001001;
DRAM[43866] = 8'b10001000;
DRAM[43867] = 8'b10001001;
DRAM[43868] = 8'b10001101;
DRAM[43869] = 8'b10010011;
DRAM[43870] = 8'b10011001;
DRAM[43871] = 8'b10011101;
DRAM[43872] = 8'b10011100;
DRAM[43873] = 8'b10100001;
DRAM[43874] = 8'b10101001;
DRAM[43875] = 8'b10110001;
DRAM[43876] = 8'b10110101;
DRAM[43877] = 8'b10110100;
DRAM[43878] = 8'b10110010;
DRAM[43879] = 8'b10110010;
DRAM[43880] = 8'b10101001;
DRAM[43881] = 8'b10101010;
DRAM[43882] = 8'b10101010;
DRAM[43883] = 8'b10101101;
DRAM[43884] = 8'b10110111;
DRAM[43885] = 8'b11000100;
DRAM[43886] = 8'b11000111;
DRAM[43887] = 8'b11000010;
DRAM[43888] = 8'b11001010;
DRAM[43889] = 8'b11010000;
DRAM[43890] = 8'b11010000;
DRAM[43891] = 8'b11000110;
DRAM[43892] = 8'b10111100;
DRAM[43893] = 8'b10110110;
DRAM[43894] = 8'b10110101;
DRAM[43895] = 8'b10110011;
DRAM[43896] = 8'b10101111;
DRAM[43897] = 8'b10100111;
DRAM[43898] = 8'b10100010;
DRAM[43899] = 8'b10100101;
DRAM[43900] = 8'b10100110;
DRAM[43901] = 8'b10100001;
DRAM[43902] = 8'b10011001;
DRAM[43903] = 8'b10010100;
DRAM[43904] = 8'b1111100;
DRAM[43905] = 8'b1111110;
DRAM[43906] = 8'b1110001;
DRAM[43907] = 8'b1011010;
DRAM[43908] = 8'b1001100;
DRAM[43909] = 8'b1001101;
DRAM[43910] = 8'b1001010;
DRAM[43911] = 8'b1000001;
DRAM[43912] = 8'b110010;
DRAM[43913] = 8'b11111;
DRAM[43914] = 8'b1101;
DRAM[43915] = 8'b110;
DRAM[43916] = 8'b110;
DRAM[43917] = 8'b100;
DRAM[43918] = 8'b1;
DRAM[43919] = 8'b0;
DRAM[43920] = 8'b0;
DRAM[43921] = 8'b0;
DRAM[43922] = 8'b0;
DRAM[43923] = 8'b0;
DRAM[43924] = 8'b0;
DRAM[43925] = 8'b0;
DRAM[43926] = 8'b0;
DRAM[43927] = 8'b0;
DRAM[43928] = 8'b1;
DRAM[43929] = 8'b0;
DRAM[43930] = 8'b0;
DRAM[43931] = 8'b0;
DRAM[43932] = 8'b10;
DRAM[43933] = 8'b1000;
DRAM[43934] = 8'b1111;
DRAM[43935] = 8'b10011;
DRAM[43936] = 8'b110001;
DRAM[43937] = 8'b1000010;
DRAM[43938] = 8'b1001110;
DRAM[43939] = 8'b1011010;
DRAM[43940] = 8'b1101100;
DRAM[43941] = 8'b1110110;
DRAM[43942] = 8'b1111101;
DRAM[43943] = 8'b10001011;
DRAM[43944] = 8'b10010111;
DRAM[43945] = 8'b10010110;
DRAM[43946] = 8'b10011110;
DRAM[43947] = 8'b10101100;
DRAM[43948] = 8'b10110101;
DRAM[43949] = 8'b10111000;
DRAM[43950] = 8'b10111111;
DRAM[43951] = 8'b11001000;
DRAM[43952] = 8'b11010100;
DRAM[43953] = 8'b11011110;
DRAM[43954] = 8'b11100011;
DRAM[43955] = 8'b11100010;
DRAM[43956] = 8'b11011110;
DRAM[43957] = 8'b11011011;
DRAM[43958] = 8'b11011110;
DRAM[43959] = 8'b11100111;
DRAM[43960] = 8'b11010001;
DRAM[43961] = 8'b10011100;
DRAM[43962] = 8'b10100100;
DRAM[43963] = 8'b10110100;
DRAM[43964] = 8'b11000011;
DRAM[43965] = 8'b11011011;
DRAM[43966] = 8'b11011110;
DRAM[43967] = 8'b11101100;
DRAM[43968] = 8'b11011001;
DRAM[43969] = 8'b11010011;
DRAM[43970] = 8'b11001101;
DRAM[43971] = 8'b11001101;
DRAM[43972] = 8'b11001111;
DRAM[43973] = 8'b11001111;
DRAM[43974] = 8'b11001011;
DRAM[43975] = 8'b11000111;
DRAM[43976] = 8'b10101010;
DRAM[43977] = 8'b10101000;
DRAM[43978] = 8'b10101110;
DRAM[43979] = 8'b10110011;
DRAM[43980] = 8'b10100111;
DRAM[43981] = 8'b10010110;
DRAM[43982] = 8'b10011011;
DRAM[43983] = 8'b10101110;
DRAM[43984] = 8'b10100110;
DRAM[43985] = 8'b10100000;
DRAM[43986] = 8'b10011011;
DRAM[43987] = 8'b10011001;
DRAM[43988] = 8'b10010101;
DRAM[43989] = 8'b10001111;
DRAM[43990] = 8'b10001101;
DRAM[43991] = 8'b10001110;
DRAM[43992] = 8'b10001111;
DRAM[43993] = 8'b10001110;
DRAM[43994] = 8'b10001100;
DRAM[43995] = 8'b10001100;
DRAM[43996] = 8'b10001101;
DRAM[43997] = 8'b10001100;
DRAM[43998] = 8'b10001001;
DRAM[43999] = 8'b10000111;
DRAM[44000] = 8'b10000111;
DRAM[44001] = 8'b10000100;
DRAM[44002] = 8'b10000010;
DRAM[44003] = 8'b10000000;
DRAM[44004] = 8'b1111111;
DRAM[44005] = 8'b1111110;
DRAM[44006] = 8'b1111011;
DRAM[44007] = 8'b1111000;
DRAM[44008] = 8'b1111010;
DRAM[44009] = 8'b1111010;
DRAM[44010] = 8'b1111011;
DRAM[44011] = 8'b1111100;
DRAM[44012] = 8'b1111110;
DRAM[44013] = 8'b10000000;
DRAM[44014] = 8'b10000010;
DRAM[44015] = 8'b10000011;
DRAM[44016] = 8'b10000010;
DRAM[44017] = 8'b10000010;
DRAM[44018] = 8'b10000100;
DRAM[44019] = 8'b10000101;
DRAM[44020] = 8'b10000110;
DRAM[44021] = 8'b10000110;
DRAM[44022] = 8'b10000110;
DRAM[44023] = 8'b10000110;
DRAM[44024] = 8'b10000110;
DRAM[44025] = 8'b10000110;
DRAM[44026] = 8'b10000110;
DRAM[44027] = 8'b10000110;
DRAM[44028] = 8'b10000111;
DRAM[44029] = 8'b10000111;
DRAM[44030] = 8'b10000111;
DRAM[44031] = 8'b10000111;
DRAM[44032] = 8'b10010011;
DRAM[44033] = 8'b10010011;
DRAM[44034] = 8'b10010011;
DRAM[44035] = 8'b10010011;
DRAM[44036] = 8'b10010100;
DRAM[44037] = 8'b10010100;
DRAM[44038] = 8'b10010100;
DRAM[44039] = 8'b10010101;
DRAM[44040] = 8'b10010101;
DRAM[44041] = 8'b10010101;
DRAM[44042] = 8'b10010111;
DRAM[44043] = 8'b10011000;
DRAM[44044] = 8'b10011001;
DRAM[44045] = 8'b10011001;
DRAM[44046] = 8'b10011001;
DRAM[44047] = 8'b10011001;
DRAM[44048] = 8'b10011011;
DRAM[44049] = 8'b10011100;
DRAM[44050] = 8'b10011100;
DRAM[44051] = 8'b10011101;
DRAM[44052] = 8'b10011110;
DRAM[44053] = 8'b10011111;
DRAM[44054] = 8'b10100000;
DRAM[44055] = 8'b10100000;
DRAM[44056] = 8'b10100001;
DRAM[44057] = 8'b10100000;
DRAM[44058] = 8'b10100000;
DRAM[44059] = 8'b10100001;
DRAM[44060] = 8'b10100001;
DRAM[44061] = 8'b10100011;
DRAM[44062] = 8'b10100100;
DRAM[44063] = 8'b10100101;
DRAM[44064] = 8'b10101000;
DRAM[44065] = 8'b10101010;
DRAM[44066] = 8'b10101110;
DRAM[44067] = 8'b10110101;
DRAM[44068] = 8'b11000010;
DRAM[44069] = 8'b11011000;
DRAM[44070] = 8'b11101111;
DRAM[44071] = 8'b11111111;
DRAM[44072] = 8'b11111101;
DRAM[44073] = 8'b11111101;
DRAM[44074] = 8'b11111101;
DRAM[44075] = 8'b11111110;
DRAM[44076] = 8'b11111110;
DRAM[44077] = 8'b11111111;
DRAM[44078] = 8'b11111111;
DRAM[44079] = 8'b11111111;
DRAM[44080] = 8'b11111110;
DRAM[44081] = 8'b11111110;
DRAM[44082] = 8'b11111110;
DRAM[44083] = 8'b11111110;
DRAM[44084] = 8'b11111110;
DRAM[44085] = 8'b11111110;
DRAM[44086] = 8'b11111110;
DRAM[44087] = 8'b11111110;
DRAM[44088] = 8'b11111100;
DRAM[44089] = 8'b11111001;
DRAM[44090] = 8'b11110110;
DRAM[44091] = 8'b11110101;
DRAM[44092] = 8'b11110100;
DRAM[44093] = 8'b11110010;
DRAM[44094] = 8'b11101101;
DRAM[44095] = 8'b11101010;
DRAM[44096] = 8'b11011110;
DRAM[44097] = 8'b11011110;
DRAM[44098] = 8'b11011111;
DRAM[44099] = 8'b11011111;
DRAM[44100] = 8'b11011101;
DRAM[44101] = 8'b11010111;
DRAM[44102] = 8'b11001111;
DRAM[44103] = 8'b11001000;
DRAM[44104] = 8'b10111011;
DRAM[44105] = 8'b10111100;
DRAM[44106] = 8'b10111100;
DRAM[44107] = 8'b10111000;
DRAM[44108] = 8'b10110011;
DRAM[44109] = 8'b10101111;
DRAM[44110] = 8'b10101101;
DRAM[44111] = 8'b10101011;
DRAM[44112] = 8'b10101111;
DRAM[44113] = 8'b10101000;
DRAM[44114] = 8'b10100000;
DRAM[44115] = 8'b10011011;
DRAM[44116] = 8'b10011001;
DRAM[44117] = 8'b10010111;
DRAM[44118] = 8'b10010011;
DRAM[44119] = 8'b10001110;
DRAM[44120] = 8'b10000101;
DRAM[44121] = 8'b10000111;
DRAM[44122] = 8'b10001000;
DRAM[44123] = 8'b10001000;
DRAM[44124] = 8'b10001001;
DRAM[44125] = 8'b10001101;
DRAM[44126] = 8'b10010110;
DRAM[44127] = 8'b10011101;
DRAM[44128] = 8'b10010111;
DRAM[44129] = 8'b10011110;
DRAM[44130] = 8'b10100110;
DRAM[44131] = 8'b10101101;
DRAM[44132] = 8'b10110010;
DRAM[44133] = 8'b10110011;
DRAM[44134] = 8'b10101111;
DRAM[44135] = 8'b10101011;
DRAM[44136] = 8'b10101101;
DRAM[44137] = 8'b10101111;
DRAM[44138] = 8'b10110010;
DRAM[44139] = 8'b10110111;
DRAM[44140] = 8'b10111110;
DRAM[44141] = 8'b11000110;
DRAM[44142] = 8'b11001001;
DRAM[44143] = 8'b11000111;
DRAM[44144] = 8'b10110111;
DRAM[44145] = 8'b11000100;
DRAM[44146] = 8'b11001011;
DRAM[44147] = 8'b11000011;
DRAM[44148] = 8'b10111000;
DRAM[44149] = 8'b10110101;
DRAM[44150] = 8'b10111011;
DRAM[44151] = 8'b11000001;
DRAM[44152] = 8'b10101001;
DRAM[44153] = 8'b10100011;
DRAM[44154] = 8'b10100000;
DRAM[44155] = 8'b10100011;
DRAM[44156] = 8'b10100100;
DRAM[44157] = 8'b10011101;
DRAM[44158] = 8'b10010101;
DRAM[44159] = 8'b10010001;
DRAM[44160] = 8'b10000101;
DRAM[44161] = 8'b10000101;
DRAM[44162] = 8'b1110111;
DRAM[44163] = 8'b1100000;
DRAM[44164] = 8'b1010100;
DRAM[44165] = 8'b1010011;
DRAM[44166] = 8'b1001011;
DRAM[44167] = 8'b111111;
DRAM[44168] = 8'b110000;
DRAM[44169] = 8'b100011;
DRAM[44170] = 8'b10100;
DRAM[44171] = 8'b1011;
DRAM[44172] = 8'b100;
DRAM[44173] = 8'b0;
DRAM[44174] = 8'b0;
DRAM[44175] = 8'b10;
DRAM[44176] = 8'b0;
DRAM[44177] = 8'b0;
DRAM[44178] = 8'b0;
DRAM[44179] = 8'b0;
DRAM[44180] = 8'b0;
DRAM[44181] = 8'b0;
DRAM[44182] = 8'b0;
DRAM[44183] = 8'b0;
DRAM[44184] = 8'b1;
DRAM[44185] = 8'b0;
DRAM[44186] = 8'b0;
DRAM[44187] = 8'b0;
DRAM[44188] = 8'b100;
DRAM[44189] = 8'b1011;
DRAM[44190] = 8'b10011;
DRAM[44191] = 8'b10111;
DRAM[44192] = 8'b110001;
DRAM[44193] = 8'b1000001;
DRAM[44194] = 8'b1001101;
DRAM[44195] = 8'b1011010;
DRAM[44196] = 8'b1101101;
DRAM[44197] = 8'b1110110;
DRAM[44198] = 8'b1111100;
DRAM[44199] = 8'b10001000;
DRAM[44200] = 8'b10000110;
DRAM[44201] = 8'b10001001;
DRAM[44202] = 8'b10010101;
DRAM[44203] = 8'b10100111;
DRAM[44204] = 8'b10101110;
DRAM[44205] = 8'b10110001;
DRAM[44206] = 8'b10111110;
DRAM[44207] = 8'b11001111;
DRAM[44208] = 8'b11010111;
DRAM[44209] = 8'b11100001;
DRAM[44210] = 8'b11100100;
DRAM[44211] = 8'b11011001;
DRAM[44212] = 8'b11010111;
DRAM[44213] = 8'b11100011;
DRAM[44214] = 8'b11100010;
DRAM[44215] = 8'b11010010;
DRAM[44216] = 8'b11010010;
DRAM[44217] = 8'b10110110;
DRAM[44218] = 8'b10111111;
DRAM[44219] = 8'b10110100;
DRAM[44220] = 8'b10111101;
DRAM[44221] = 8'b11101001;
DRAM[44222] = 8'b11101001;
DRAM[44223] = 8'b11011111;
DRAM[44224] = 8'b11100010;
DRAM[44225] = 8'b11100011;
DRAM[44226] = 8'b11011110;
DRAM[44227] = 8'b11010000;
DRAM[44228] = 8'b11000010;
DRAM[44229] = 8'b10111110;
DRAM[44230] = 8'b11000101;
DRAM[44231] = 8'b11001101;
DRAM[44232] = 8'b11000011;
DRAM[44233] = 8'b10101010;
DRAM[44234] = 8'b10011100;
DRAM[44235] = 8'b10100100;
DRAM[44236] = 8'b10101001;
DRAM[44237] = 8'b10100001;
DRAM[44238] = 8'b10100001;
DRAM[44239] = 8'b10101011;
DRAM[44240] = 8'b10100011;
DRAM[44241] = 8'b10011111;
DRAM[44242] = 8'b10011101;
DRAM[44243] = 8'b10011100;
DRAM[44244] = 8'b10010111;
DRAM[44245] = 8'b10001111;
DRAM[44246] = 8'b10001010;
DRAM[44247] = 8'b10001011;
DRAM[44248] = 8'b10001110;
DRAM[44249] = 8'b10001100;
DRAM[44250] = 8'b10001011;
DRAM[44251] = 8'b10001011;
DRAM[44252] = 8'b10001011;
DRAM[44253] = 8'b10001010;
DRAM[44254] = 8'b10001000;
DRAM[44255] = 8'b10000101;
DRAM[44256] = 8'b10000111;
DRAM[44257] = 8'b10000101;
DRAM[44258] = 8'b10000010;
DRAM[44259] = 8'b10000001;
DRAM[44260] = 8'b10000000;
DRAM[44261] = 8'b1111111;
DRAM[44262] = 8'b1111100;
DRAM[44263] = 8'b1111010;
DRAM[44264] = 8'b1111101;
DRAM[44265] = 8'b1111101;
DRAM[44266] = 8'b1111101;
DRAM[44267] = 8'b1111101;
DRAM[44268] = 8'b1111101;
DRAM[44269] = 8'b1111111;
DRAM[44270] = 8'b10000000;
DRAM[44271] = 8'b10000001;
DRAM[44272] = 8'b10000011;
DRAM[44273] = 8'b10000011;
DRAM[44274] = 8'b10000101;
DRAM[44275] = 8'b10000110;
DRAM[44276] = 8'b10000110;
DRAM[44277] = 8'b10000111;
DRAM[44278] = 8'b10000110;
DRAM[44279] = 8'b10000110;
DRAM[44280] = 8'b10000110;
DRAM[44281] = 8'b10000110;
DRAM[44282] = 8'b10000111;
DRAM[44283] = 8'b10000111;
DRAM[44284] = 8'b10001000;
DRAM[44285] = 8'b10001000;
DRAM[44286] = 8'b10001001;
DRAM[44287] = 8'b10001001;
DRAM[44288] = 8'b10010010;
DRAM[44289] = 8'b10010010;
DRAM[44290] = 8'b10010010;
DRAM[44291] = 8'b10010011;
DRAM[44292] = 8'b10010011;
DRAM[44293] = 8'b10010011;
DRAM[44294] = 8'b10010100;
DRAM[44295] = 8'b10010100;
DRAM[44296] = 8'b10010100;
DRAM[44297] = 8'b10010101;
DRAM[44298] = 8'b10010111;
DRAM[44299] = 8'b10011000;
DRAM[44300] = 8'b10011001;
DRAM[44301] = 8'b10011001;
DRAM[44302] = 8'b10011001;
DRAM[44303] = 8'b10011001;
DRAM[44304] = 8'b10011010;
DRAM[44305] = 8'b10011010;
DRAM[44306] = 8'b10011011;
DRAM[44307] = 8'b10011100;
DRAM[44308] = 8'b10011101;
DRAM[44309] = 8'b10011110;
DRAM[44310] = 8'b10011111;
DRAM[44311] = 8'b10100000;
DRAM[44312] = 8'b10100000;
DRAM[44313] = 8'b10100000;
DRAM[44314] = 8'b10100000;
DRAM[44315] = 8'b10100000;
DRAM[44316] = 8'b10100001;
DRAM[44317] = 8'b10100010;
DRAM[44318] = 8'b10100100;
DRAM[44319] = 8'b10100100;
DRAM[44320] = 8'b10101001;
DRAM[44321] = 8'b10101100;
DRAM[44322] = 8'b10110001;
DRAM[44323] = 8'b10111001;
DRAM[44324] = 8'b11000110;
DRAM[44325] = 8'b11011010;
DRAM[44326] = 8'b11110000;
DRAM[44327] = 8'b11111110;
DRAM[44328] = 8'b11111101;
DRAM[44329] = 8'b11111101;
DRAM[44330] = 8'b11111101;
DRAM[44331] = 8'b11111110;
DRAM[44332] = 8'b11111110;
DRAM[44333] = 8'b11111111;
DRAM[44334] = 8'b11111111;
DRAM[44335] = 8'b11111111;
DRAM[44336] = 8'b11111111;
DRAM[44337] = 8'b11111111;
DRAM[44338] = 8'b11111110;
DRAM[44339] = 8'b11111110;
DRAM[44340] = 8'b11111110;
DRAM[44341] = 8'b11111110;
DRAM[44342] = 8'b11111101;
DRAM[44343] = 8'b11111101;
DRAM[44344] = 8'b11111100;
DRAM[44345] = 8'b11111000;
DRAM[44346] = 8'b11110100;
DRAM[44347] = 8'b11110011;
DRAM[44348] = 8'b11110100;
DRAM[44349] = 8'b11110011;
DRAM[44350] = 8'b11101101;
DRAM[44351] = 8'b11101000;
DRAM[44352] = 8'b11100111;
DRAM[44353] = 8'b11100100;
DRAM[44354] = 8'b11100000;
DRAM[44355] = 8'b11011101;
DRAM[44356] = 8'b11011000;
DRAM[44357] = 8'b11010010;
DRAM[44358] = 8'b11001011;
DRAM[44359] = 8'b11000110;
DRAM[44360] = 8'b10111011;
DRAM[44361] = 8'b10111100;
DRAM[44362] = 8'b10111010;
DRAM[44363] = 8'b10110110;
DRAM[44364] = 8'b10110101;
DRAM[44365] = 8'b10110110;
DRAM[44366] = 8'b10110101;
DRAM[44367] = 8'b10110001;
DRAM[44368] = 8'b10100101;
DRAM[44369] = 8'b10100010;
DRAM[44370] = 8'b10011111;
DRAM[44371] = 8'b10100000;
DRAM[44372] = 8'b10100000;
DRAM[44373] = 8'b10011010;
DRAM[44374] = 8'b10001110;
DRAM[44375] = 8'b10000100;
DRAM[44376] = 8'b10001100;
DRAM[44377] = 8'b10001110;
DRAM[44378] = 8'b10001110;
DRAM[44379] = 8'b10001011;
DRAM[44380] = 8'b10000111;
DRAM[44381] = 8'b10000111;
DRAM[44382] = 8'b10001101;
DRAM[44383] = 8'b10010010;
DRAM[44384] = 8'b10010000;
DRAM[44385] = 8'b10010110;
DRAM[44386] = 8'b10011101;
DRAM[44387] = 8'b10100010;
DRAM[44388] = 8'b10100111;
DRAM[44389] = 8'b10101010;
DRAM[44390] = 8'b10100110;
DRAM[44391] = 8'b10100000;
DRAM[44392] = 8'b10101011;
DRAM[44393] = 8'b10101010;
DRAM[44394] = 8'b10101011;
DRAM[44395] = 8'b10110001;
DRAM[44396] = 8'b10111010;
DRAM[44397] = 8'b11000001;
DRAM[44398] = 8'b11000011;
DRAM[44399] = 8'b11000001;
DRAM[44400] = 8'b10110110;
DRAM[44401] = 8'b11000101;
DRAM[44402] = 8'b11010000;
DRAM[44403] = 8'b11001011;
DRAM[44404] = 8'b10111110;
DRAM[44405] = 8'b10110101;
DRAM[44406] = 8'b10110011;
DRAM[44407] = 8'b10110011;
DRAM[44408] = 8'b10101000;
DRAM[44409] = 8'b10100001;
DRAM[44410] = 8'b10011101;
DRAM[44411] = 8'b10011111;
DRAM[44412] = 8'b10011110;
DRAM[44413] = 8'b10010111;
DRAM[44414] = 8'b10010001;
DRAM[44415] = 8'b10001111;
DRAM[44416] = 8'b10001011;
DRAM[44417] = 8'b1111101;
DRAM[44418] = 8'b1110100;
DRAM[44419] = 8'b1110010;
DRAM[44420] = 8'b1100111;
DRAM[44421] = 8'b1001111;
DRAM[44422] = 8'b1000000;
DRAM[44423] = 8'b111110;
DRAM[44424] = 8'b101110;
DRAM[44425] = 8'b100100;
DRAM[44426] = 8'b11001;
DRAM[44427] = 8'b1111;
DRAM[44428] = 8'b101;
DRAM[44429] = 8'b0;
DRAM[44430] = 8'b0;
DRAM[44431] = 8'b11;
DRAM[44432] = 8'b0;
DRAM[44433] = 8'b0;
DRAM[44434] = 8'b0;
DRAM[44435] = 8'b0;
DRAM[44436] = 8'b0;
DRAM[44437] = 8'b0;
DRAM[44438] = 8'b0;
DRAM[44439] = 8'b0;
DRAM[44440] = 8'b0;
DRAM[44441] = 8'b0;
DRAM[44442] = 8'b0;
DRAM[44443] = 8'b1;
DRAM[44444] = 8'b101;
DRAM[44445] = 8'b1101;
DRAM[44446] = 8'b10100;
DRAM[44447] = 8'b11001;
DRAM[44448] = 8'b101011;
DRAM[44449] = 8'b111010;
DRAM[44450] = 8'b1000101;
DRAM[44451] = 8'b1010000;
DRAM[44452] = 8'b1100001;
DRAM[44453] = 8'b1101000;
DRAM[44454] = 8'b1101110;
DRAM[44455] = 8'b1111010;
DRAM[44456] = 8'b1111000;
DRAM[44457] = 8'b10000001;
DRAM[44458] = 8'b10010100;
DRAM[44459] = 8'b10100110;
DRAM[44460] = 8'b10101100;
DRAM[44461] = 8'b10101110;
DRAM[44462] = 8'b10111001;
DRAM[44463] = 8'b11001000;
DRAM[44464] = 8'b11011100;
DRAM[44465] = 8'b11100011;
DRAM[44466] = 8'b11100100;
DRAM[44467] = 8'b11010110;
DRAM[44468] = 8'b11010001;
DRAM[44469] = 8'b11100010;
DRAM[44470] = 8'b11011101;
DRAM[44471] = 8'b10111101;
DRAM[44472] = 8'b10110011;
DRAM[44473] = 8'b10110110;
DRAM[44474] = 8'b11010000;
DRAM[44475] = 8'b11011101;
DRAM[44476] = 8'b11100001;
DRAM[44477] = 8'b11101000;
DRAM[44478] = 8'b11100001;
DRAM[44479] = 8'b11011111;
DRAM[44480] = 8'b11100110;
DRAM[44481] = 8'b11011001;
DRAM[44482] = 8'b11001011;
DRAM[44483] = 8'b11000111;
DRAM[44484] = 8'b11001110;
DRAM[44485] = 8'b11001110;
DRAM[44486] = 8'b10111111;
DRAM[44487] = 8'b10101100;
DRAM[44488] = 8'b10111010;
DRAM[44489] = 8'b10110101;
DRAM[44490] = 8'b10101100;
DRAM[44491] = 8'b10100011;
DRAM[44492] = 8'b10100010;
DRAM[44493] = 8'b10100110;
DRAM[44494] = 8'b10100110;
DRAM[44495] = 8'b10100010;
DRAM[44496] = 8'b10011100;
DRAM[44497] = 8'b10011011;
DRAM[44498] = 8'b10011100;
DRAM[44499] = 8'b10011101;
DRAM[44500] = 8'b10011000;
DRAM[44501] = 8'b10010000;
DRAM[44502] = 8'b10001101;
DRAM[44503] = 8'b10001111;
DRAM[44504] = 8'b10001101;
DRAM[44505] = 8'b10001011;
DRAM[44506] = 8'b10001010;
DRAM[44507] = 8'b10001010;
DRAM[44508] = 8'b10001010;
DRAM[44509] = 8'b10001001;
DRAM[44510] = 8'b10000111;
DRAM[44511] = 8'b10000100;
DRAM[44512] = 8'b10000110;
DRAM[44513] = 8'b10000100;
DRAM[44514] = 8'b10000001;
DRAM[44515] = 8'b10000001;
DRAM[44516] = 8'b10000001;
DRAM[44517] = 8'b10000000;
DRAM[44518] = 8'b1111110;
DRAM[44519] = 8'b1111011;
DRAM[44520] = 8'b1111111;
DRAM[44521] = 8'b1111110;
DRAM[44522] = 8'b1111101;
DRAM[44523] = 8'b1111101;
DRAM[44524] = 8'b1111101;
DRAM[44525] = 8'b1111110;
DRAM[44526] = 8'b10000000;
DRAM[44527] = 8'b10000001;
DRAM[44528] = 8'b10000100;
DRAM[44529] = 8'b10000100;
DRAM[44530] = 8'b10000101;
DRAM[44531] = 8'b10000110;
DRAM[44532] = 8'b10000111;
DRAM[44533] = 8'b10000111;
DRAM[44534] = 8'b10000110;
DRAM[44535] = 8'b10000110;
DRAM[44536] = 8'b10000110;
DRAM[44537] = 8'b10000111;
DRAM[44538] = 8'b10000111;
DRAM[44539] = 8'b10001000;
DRAM[44540] = 8'b10001001;
DRAM[44541] = 8'b10001001;
DRAM[44542] = 8'b10001010;
DRAM[44543] = 8'b10001010;
DRAM[44544] = 8'b10010001;
DRAM[44545] = 8'b10010001;
DRAM[44546] = 8'b10010010;
DRAM[44547] = 8'b10010010;
DRAM[44548] = 8'b10010010;
DRAM[44549] = 8'b10010011;
DRAM[44550] = 8'b10010011;
DRAM[44551] = 8'b10010011;
DRAM[44552] = 8'b10010101;
DRAM[44553] = 8'b10010110;
DRAM[44554] = 8'b10010111;
DRAM[44555] = 8'b10011000;
DRAM[44556] = 8'b10011001;
DRAM[44557] = 8'b10011001;
DRAM[44558] = 8'b10011001;
DRAM[44559] = 8'b10011001;
DRAM[44560] = 8'b10011001;
DRAM[44561] = 8'b10011001;
DRAM[44562] = 8'b10011010;
DRAM[44563] = 8'b10011100;
DRAM[44564] = 8'b10011101;
DRAM[44565] = 8'b10011110;
DRAM[44566] = 8'b10011111;
DRAM[44567] = 8'b10100000;
DRAM[44568] = 8'b10100000;
DRAM[44569] = 8'b10100000;
DRAM[44570] = 8'b10100000;
DRAM[44571] = 8'b10100000;
DRAM[44572] = 8'b10100001;
DRAM[44573] = 8'b10100010;
DRAM[44574] = 8'b10100011;
DRAM[44575] = 8'b10100100;
DRAM[44576] = 8'b10101011;
DRAM[44577] = 8'b10101110;
DRAM[44578] = 8'b10110110;
DRAM[44579] = 8'b11000101;
DRAM[44580] = 8'b11011000;
DRAM[44581] = 8'b11101001;
DRAM[44582] = 8'b11110110;
DRAM[44583] = 8'b11111100;
DRAM[44584] = 8'b11111101;
DRAM[44585] = 8'b11111101;
DRAM[44586] = 8'b11111101;
DRAM[44587] = 8'b11111110;
DRAM[44588] = 8'b11111110;
DRAM[44589] = 8'b11111111;
DRAM[44590] = 8'b11111111;
DRAM[44591] = 8'b11111111;
DRAM[44592] = 8'b11111111;
DRAM[44593] = 8'b11111111;
DRAM[44594] = 8'b11111111;
DRAM[44595] = 8'b11111110;
DRAM[44596] = 8'b11111110;
DRAM[44597] = 8'b11111101;
DRAM[44598] = 8'b11111101;
DRAM[44599] = 8'b11111101;
DRAM[44600] = 8'b11111001;
DRAM[44601] = 8'b11111000;
DRAM[44602] = 8'b11110110;
DRAM[44603] = 8'b11110100;
DRAM[44604] = 8'b11110010;
DRAM[44605] = 8'b11101111;
DRAM[44606] = 8'b11101100;
DRAM[44607] = 8'b11101010;
DRAM[44608] = 8'b11101100;
DRAM[44609] = 8'b11100101;
DRAM[44610] = 8'b11011011;
DRAM[44611] = 8'b11010010;
DRAM[44612] = 8'b11001101;
DRAM[44613] = 8'b11001010;
DRAM[44614] = 8'b11001000;
DRAM[44615] = 8'b11000111;
DRAM[44616] = 8'b10111010;
DRAM[44617] = 8'b10111011;
DRAM[44618] = 8'b10110111;
DRAM[44619] = 8'b10110100;
DRAM[44620] = 8'b10110111;
DRAM[44621] = 8'b10111110;
DRAM[44622] = 8'b10111110;
DRAM[44623] = 8'b10111001;
DRAM[44624] = 8'b10100010;
DRAM[44625] = 8'b10100001;
DRAM[44626] = 8'b10100010;
DRAM[44627] = 8'b10100011;
DRAM[44628] = 8'b10100010;
DRAM[44629] = 8'b10011101;
DRAM[44630] = 8'b10010101;
DRAM[44631] = 8'b10001110;
DRAM[44632] = 8'b10010010;
DRAM[44633] = 8'b10010000;
DRAM[44634] = 8'b10001101;
DRAM[44635] = 8'b10001011;
DRAM[44636] = 8'b10001001;
DRAM[44637] = 8'b10001000;
DRAM[44638] = 8'b10001000;
DRAM[44639] = 8'b10001000;
DRAM[44640] = 8'b10010001;
DRAM[44641] = 8'b10011000;
DRAM[44642] = 8'b10011110;
DRAM[44643] = 8'b10100100;
DRAM[44644] = 8'b10101100;
DRAM[44645] = 8'b10110100;
DRAM[44646] = 8'b10110011;
DRAM[44647] = 8'b10101100;
DRAM[44648] = 8'b10011111;
DRAM[44649] = 8'b10010100;
DRAM[44650] = 8'b10001111;
DRAM[44651] = 8'b10011010;
DRAM[44652] = 8'b10101111;
DRAM[44653] = 8'b10111101;
DRAM[44654] = 8'b10111110;
DRAM[44655] = 8'b10111011;
DRAM[44656] = 8'b11000001;
DRAM[44657] = 8'b11001001;
DRAM[44658] = 8'b11001110;
DRAM[44659] = 8'b11001010;
DRAM[44660] = 8'b11000000;
DRAM[44661] = 8'b10110101;
DRAM[44662] = 8'b10101001;
DRAM[44663] = 8'b10011111;
DRAM[44664] = 8'b10100100;
DRAM[44665] = 8'b10011100;
DRAM[44666] = 8'b10010110;
DRAM[44667] = 8'b10010101;
DRAM[44668] = 8'b10010100;
DRAM[44669] = 8'b10010000;
DRAM[44670] = 8'b10001101;
DRAM[44671] = 8'b10001101;
DRAM[44672] = 8'b10000110;
DRAM[44673] = 8'b1111001;
DRAM[44674] = 8'b1110001;
DRAM[44675] = 8'b1101111;
DRAM[44676] = 8'b1100001;
DRAM[44677] = 8'b1001010;
DRAM[44678] = 8'b111110;
DRAM[44679] = 8'b111111;
DRAM[44680] = 8'b101111;
DRAM[44681] = 8'b100100;
DRAM[44682] = 8'b11001;
DRAM[44683] = 8'b10001;
DRAM[44684] = 8'b1010;
DRAM[44685] = 8'b11;
DRAM[44686] = 8'b0;
DRAM[44687] = 8'b10;
DRAM[44688] = 8'b0;
DRAM[44689] = 8'b0;
DRAM[44690] = 8'b0;
DRAM[44691] = 8'b0;
DRAM[44692] = 8'b0;
DRAM[44693] = 8'b0;
DRAM[44694] = 8'b0;
DRAM[44695] = 8'b0;
DRAM[44696] = 8'b0;
DRAM[44697] = 8'b0;
DRAM[44698] = 8'b0;
DRAM[44699] = 8'b10;
DRAM[44700] = 8'b111;
DRAM[44701] = 8'b1110;
DRAM[44702] = 8'b10100;
DRAM[44703] = 8'b11001;
DRAM[44704] = 8'b100110;
DRAM[44705] = 8'b110101;
DRAM[44706] = 8'b111110;
DRAM[44707] = 8'b1000101;
DRAM[44708] = 8'b1010011;
DRAM[44709] = 8'b1011011;
DRAM[44710] = 8'b1100100;
DRAM[44711] = 8'b1110011;
DRAM[44712] = 8'b1111000;
DRAM[44713] = 8'b10000001;
DRAM[44714] = 8'b10010000;
DRAM[44715] = 8'b10011110;
DRAM[44716] = 8'b10101000;
DRAM[44717] = 8'b10110001;
DRAM[44718] = 8'b10111011;
DRAM[44719] = 8'b11000100;
DRAM[44720] = 8'b11011001;
DRAM[44721] = 8'b11011001;
DRAM[44722] = 8'b11011111;
DRAM[44723] = 8'b11011001;
DRAM[44724] = 8'b11010000;
DRAM[44725] = 8'b11011011;
DRAM[44726] = 8'b11011000;
DRAM[44727] = 8'b10111011;
DRAM[44728] = 8'b10100101;
DRAM[44729] = 8'b10110000;
DRAM[44730] = 8'b11000010;
DRAM[44731] = 8'b11101101;
DRAM[44732] = 8'b11111100;
DRAM[44733] = 8'b11100011;
DRAM[44734] = 8'b11011111;
DRAM[44735] = 8'b11101010;
DRAM[44736] = 8'b11011100;
DRAM[44737] = 8'b11011001;
DRAM[44738] = 8'b11001100;
DRAM[44739] = 8'b10111001;
DRAM[44740] = 8'b10110000;
DRAM[44741] = 8'b10110110;
DRAM[44742] = 8'b10111111;
DRAM[44743] = 8'b11000100;
DRAM[44744] = 8'b10100110;
DRAM[44745] = 8'b10110010;
DRAM[44746] = 8'b10111010;
DRAM[44747] = 8'b10110100;
DRAM[44748] = 8'b10100110;
DRAM[44749] = 8'b10011101;
DRAM[44750] = 8'b10011101;
DRAM[44751] = 8'b10100000;
DRAM[44752] = 8'b10011100;
DRAM[44753] = 8'b10011011;
DRAM[44754] = 8'b10011011;
DRAM[44755] = 8'b10011011;
DRAM[44756] = 8'b10010110;
DRAM[44757] = 8'b10001111;
DRAM[44758] = 8'b10001110;
DRAM[44759] = 8'b10010010;
DRAM[44760] = 8'b10001100;
DRAM[44761] = 8'b10001010;
DRAM[44762] = 8'b10001001;
DRAM[44763] = 8'b10001001;
DRAM[44764] = 8'b10001001;
DRAM[44765] = 8'b10001000;
DRAM[44766] = 8'b10000110;
DRAM[44767] = 8'b10000011;
DRAM[44768] = 8'b10000011;
DRAM[44769] = 8'b10000001;
DRAM[44770] = 8'b1111111;
DRAM[44771] = 8'b1111111;
DRAM[44772] = 8'b10000000;
DRAM[44773] = 8'b1111111;
DRAM[44774] = 8'b1111110;
DRAM[44775] = 8'b1111100;
DRAM[44776] = 8'b1111110;
DRAM[44777] = 8'b1111101;
DRAM[44778] = 8'b1111100;
DRAM[44779] = 8'b1111100;
DRAM[44780] = 8'b1111101;
DRAM[44781] = 8'b10000000;
DRAM[44782] = 8'b10000010;
DRAM[44783] = 8'b10000100;
DRAM[44784] = 8'b10000100;
DRAM[44785] = 8'b10000101;
DRAM[44786] = 8'b10000110;
DRAM[44787] = 8'b10000111;
DRAM[44788] = 8'b10000111;
DRAM[44789] = 8'b10000111;
DRAM[44790] = 8'b10000110;
DRAM[44791] = 8'b10000110;
DRAM[44792] = 8'b10000110;
DRAM[44793] = 8'b10000111;
DRAM[44794] = 8'b10000111;
DRAM[44795] = 8'b10001000;
DRAM[44796] = 8'b10001001;
DRAM[44797] = 8'b10001010;
DRAM[44798] = 8'b10001011;
DRAM[44799] = 8'b10001011;
DRAM[44800] = 8'b10010001;
DRAM[44801] = 8'b10010001;
DRAM[44802] = 8'b10010001;
DRAM[44803] = 8'b10010010;
DRAM[44804] = 8'b10010010;
DRAM[44805] = 8'b10010010;
DRAM[44806] = 8'b10010011;
DRAM[44807] = 8'b10010011;
DRAM[44808] = 8'b10010101;
DRAM[44809] = 8'b10010110;
DRAM[44810] = 8'b10010111;
DRAM[44811] = 8'b10011000;
DRAM[44812] = 8'b10011001;
DRAM[44813] = 8'b10011010;
DRAM[44814] = 8'b10011001;
DRAM[44815] = 8'b10011001;
DRAM[44816] = 8'b10011000;
DRAM[44817] = 8'b10011001;
DRAM[44818] = 8'b10011010;
DRAM[44819] = 8'b10011011;
DRAM[44820] = 8'b10011101;
DRAM[44821] = 8'b10011110;
DRAM[44822] = 8'b10011111;
DRAM[44823] = 8'b10011111;
DRAM[44824] = 8'b10100000;
DRAM[44825] = 8'b10100000;
DRAM[44826] = 8'b10011111;
DRAM[44827] = 8'b10100000;
DRAM[44828] = 8'b10100001;
DRAM[44829] = 8'b10100010;
DRAM[44830] = 8'b10100011;
DRAM[44831] = 8'b10100100;
DRAM[44832] = 8'b10101101;
DRAM[44833] = 8'b10101111;
DRAM[44834] = 8'b10111010;
DRAM[44835] = 8'b11010000;
DRAM[44836] = 8'b11101001;
DRAM[44837] = 8'b11111001;
DRAM[44838] = 8'b11111100;
DRAM[44839] = 8'b11111001;
DRAM[44840] = 8'b11111101;
DRAM[44841] = 8'b11111101;
DRAM[44842] = 8'b11111101;
DRAM[44843] = 8'b11111110;
DRAM[44844] = 8'b11111110;
DRAM[44845] = 8'b11111111;
DRAM[44846] = 8'b11111111;
DRAM[44847] = 8'b11111111;
DRAM[44848] = 8'b11111111;
DRAM[44849] = 8'b11111111;
DRAM[44850] = 8'b11111111;
DRAM[44851] = 8'b11111110;
DRAM[44852] = 8'b11111110;
DRAM[44853] = 8'b11111101;
DRAM[44854] = 8'b11111101;
DRAM[44855] = 8'b11111101;
DRAM[44856] = 8'b11110110;
DRAM[44857] = 8'b11111000;
DRAM[44858] = 8'b11111001;
DRAM[44859] = 8'b11110110;
DRAM[44860] = 8'b11110000;
DRAM[44861] = 8'b11101011;
DRAM[44862] = 8'b11101011;
DRAM[44863] = 8'b11101100;
DRAM[44864] = 8'b11011100;
DRAM[44865] = 8'b11011100;
DRAM[44866] = 8'b11011010;
DRAM[44867] = 8'b11011000;
DRAM[44868] = 8'b11010011;
DRAM[44869] = 8'b11001011;
DRAM[44870] = 8'b11000001;
DRAM[44871] = 8'b10111010;
DRAM[44872] = 8'b10111110;
DRAM[44873] = 8'b10111100;
DRAM[44874] = 8'b10110100;
DRAM[44875] = 8'b10101110;
DRAM[44876] = 8'b10110000;
DRAM[44877] = 8'b10110111;
DRAM[44878] = 8'b10110101;
DRAM[44879] = 8'b10101101;
DRAM[44880] = 8'b10110000;
DRAM[44881] = 8'b10101110;
DRAM[44882] = 8'b10101010;
DRAM[44883] = 8'b10100011;
DRAM[44884] = 8'b10011100;
DRAM[44885] = 8'b10011001;
DRAM[44886] = 8'b10011001;
DRAM[44887] = 8'b10011010;
DRAM[44888] = 8'b10001100;
DRAM[44889] = 8'b10000111;
DRAM[44890] = 8'b10000011;
DRAM[44891] = 8'b10000100;
DRAM[44892] = 8'b10001000;
DRAM[44893] = 8'b10001010;
DRAM[44894] = 8'b10000111;
DRAM[44895] = 8'b10000011;
DRAM[44896] = 8'b10000011;
DRAM[44897] = 8'b10001010;
DRAM[44898] = 8'b10010001;
DRAM[44899] = 8'b10011001;
DRAM[44900] = 8'b10100101;
DRAM[44901] = 8'b10110001;
DRAM[44902] = 8'b10110100;
DRAM[44903] = 8'b10101111;
DRAM[44904] = 8'b10010101;
DRAM[44905] = 8'b10000100;
DRAM[44906] = 8'b1111010;
DRAM[44907] = 8'b10001010;
DRAM[44908] = 8'b10101010;
DRAM[44909] = 8'b11000001;
DRAM[44910] = 8'b11000100;
DRAM[44911] = 8'b10111110;
DRAM[44912] = 8'b11000010;
DRAM[44913] = 8'b11000010;
DRAM[44914] = 8'b11000000;
DRAM[44915] = 8'b10111101;
DRAM[44916] = 8'b10111101;
DRAM[44917] = 8'b10111010;
DRAM[44918] = 8'b10101101;
DRAM[44919] = 8'b10100000;
DRAM[44920] = 8'b10011100;
DRAM[44921] = 8'b10010100;
DRAM[44922] = 8'b10001101;
DRAM[44923] = 8'b10001100;
DRAM[44924] = 8'b10001100;
DRAM[44925] = 8'b10001010;
DRAM[44926] = 8'b10001011;
DRAM[44927] = 8'b10001110;
DRAM[44928] = 8'b1111111;
DRAM[44929] = 8'b10000010;
DRAM[44930] = 8'b1110111;
DRAM[44931] = 8'b1011111;
DRAM[44932] = 8'b1001111;
DRAM[44933] = 8'b1001110;
DRAM[44934] = 8'b1001011;
DRAM[44935] = 8'b1000011;
DRAM[44936] = 8'b110001;
DRAM[44937] = 8'b100100;
DRAM[44938] = 8'b10111;
DRAM[44939] = 8'b10010;
DRAM[44940] = 8'b1111;
DRAM[44941] = 8'b1001;
DRAM[44942] = 8'b11;
DRAM[44943] = 8'b0;
DRAM[44944] = 8'b0;
DRAM[44945] = 8'b0;
DRAM[44946] = 8'b0;
DRAM[44947] = 8'b0;
DRAM[44948] = 8'b0;
DRAM[44949] = 8'b0;
DRAM[44950] = 8'b0;
DRAM[44951] = 8'b0;
DRAM[44952] = 8'b0;
DRAM[44953] = 8'b0;
DRAM[44954] = 8'b0;
DRAM[44955] = 8'b10;
DRAM[44956] = 8'b111;
DRAM[44957] = 8'b1110;
DRAM[44958] = 8'b10100;
DRAM[44959] = 8'b11000;
DRAM[44960] = 8'b100101;
DRAM[44961] = 8'b110011;
DRAM[44962] = 8'b111010;
DRAM[44963] = 8'b1000000;
DRAM[44964] = 8'b1001101;
DRAM[44965] = 8'b1010111;
DRAM[44966] = 8'b1100100;
DRAM[44967] = 8'b1110111;
DRAM[44968] = 8'b10000000;
DRAM[44969] = 8'b10000100;
DRAM[44970] = 8'b10001011;
DRAM[44971] = 8'b10010011;
DRAM[44972] = 8'b10100010;
DRAM[44973] = 8'b10110101;
DRAM[44974] = 8'b11000011;
DRAM[44975] = 8'b11001001;
DRAM[44976] = 8'b11010010;
DRAM[44977] = 8'b11001100;
DRAM[44978] = 8'b11011001;
DRAM[44979] = 8'b11011110;
DRAM[44980] = 8'b11010011;
DRAM[44981] = 8'b11010111;
DRAM[44982] = 8'b11011000;
DRAM[44983] = 8'b11000100;
DRAM[44984] = 8'b10110111;
DRAM[44985] = 8'b11001100;
DRAM[44986] = 8'b10110100;
DRAM[44987] = 8'b11000001;
DRAM[44988] = 8'b11100000;
DRAM[44989] = 8'b11100110;
DRAM[44990] = 8'b11110011;
DRAM[44991] = 8'b11101101;
DRAM[44992] = 8'b11011000;
DRAM[44993] = 8'b11011111;
DRAM[44994] = 8'b11011101;
DRAM[44995] = 8'b11001110;
DRAM[44996] = 8'b10111101;
DRAM[44997] = 8'b10110100;
DRAM[44998] = 8'b10101111;
DRAM[44999] = 8'b10101011;
DRAM[45000] = 8'b10101110;
DRAM[45001] = 8'b10011111;
DRAM[45002] = 8'b10100000;
DRAM[45003] = 8'b10110010;
DRAM[45004] = 8'b10110010;
DRAM[45005] = 8'b10100000;
DRAM[45006] = 8'b10011101;
DRAM[45007] = 8'b10101011;
DRAM[45008] = 8'b10100010;
DRAM[45009] = 8'b10011110;
DRAM[45010] = 8'b10011100;
DRAM[45011] = 8'b10011001;
DRAM[45012] = 8'b10010010;
DRAM[45013] = 8'b10001011;
DRAM[45014] = 8'b10001100;
DRAM[45015] = 8'b10010010;
DRAM[45016] = 8'b10001011;
DRAM[45017] = 8'b10001010;
DRAM[45018] = 8'b10001001;
DRAM[45019] = 8'b10001001;
DRAM[45020] = 8'b10001001;
DRAM[45021] = 8'b10001000;
DRAM[45022] = 8'b10000101;
DRAM[45023] = 8'b10000011;
DRAM[45024] = 8'b10000000;
DRAM[45025] = 8'b1111111;
DRAM[45026] = 8'b1111101;
DRAM[45027] = 8'b1111101;
DRAM[45028] = 8'b1111110;
DRAM[45029] = 8'b1111111;
DRAM[45030] = 8'b1111101;
DRAM[45031] = 8'b1111100;
DRAM[45032] = 8'b1111100;
DRAM[45033] = 8'b1111100;
DRAM[45034] = 8'b1111011;
DRAM[45035] = 8'b1111100;
DRAM[45036] = 8'b1111110;
DRAM[45037] = 8'b10000001;
DRAM[45038] = 8'b10000100;
DRAM[45039] = 8'b10000110;
DRAM[45040] = 8'b10000101;
DRAM[45041] = 8'b10000101;
DRAM[45042] = 8'b10000110;
DRAM[45043] = 8'b10000111;
DRAM[45044] = 8'b10000111;
DRAM[45045] = 8'b10000111;
DRAM[45046] = 8'b10000110;
DRAM[45047] = 8'b10000110;
DRAM[45048] = 8'b10000111;
DRAM[45049] = 8'b10000111;
DRAM[45050] = 8'b10001000;
DRAM[45051] = 8'b10001001;
DRAM[45052] = 8'b10001010;
DRAM[45053] = 8'b10001010;
DRAM[45054] = 8'b10001011;
DRAM[45055] = 8'b10001100;
DRAM[45056] = 8'b10010001;
DRAM[45057] = 8'b10010000;
DRAM[45058] = 8'b10010000;
DRAM[45059] = 8'b10010000;
DRAM[45060] = 8'b10010000;
DRAM[45061] = 8'b10010001;
DRAM[45062] = 8'b10010010;
DRAM[45063] = 8'b10010011;
DRAM[45064] = 8'b10010100;
DRAM[45065] = 8'b10010100;
DRAM[45066] = 8'b10010110;
DRAM[45067] = 8'b10010111;
DRAM[45068] = 8'b10011000;
DRAM[45069] = 8'b10011001;
DRAM[45070] = 8'b10011001;
DRAM[45071] = 8'b10011001;
DRAM[45072] = 8'b10011000;
DRAM[45073] = 8'b10011000;
DRAM[45074] = 8'b10011001;
DRAM[45075] = 8'b10011010;
DRAM[45076] = 8'b10011011;
DRAM[45077] = 8'b10011011;
DRAM[45078] = 8'b10011100;
DRAM[45079] = 8'b10011100;
DRAM[45080] = 8'b10011111;
DRAM[45081] = 8'b10011101;
DRAM[45082] = 8'b10011100;
DRAM[45083] = 8'b10011110;
DRAM[45084] = 8'b10100010;
DRAM[45085] = 8'b10100011;
DRAM[45086] = 8'b10100001;
DRAM[45087] = 8'b10011110;
DRAM[45088] = 8'b10100001;
DRAM[45089] = 8'b10100011;
DRAM[45090] = 8'b10110100;
DRAM[45091] = 8'b11010011;
DRAM[45092] = 8'b11101110;
DRAM[45093] = 8'b11111001;
DRAM[45094] = 8'b11111011;
DRAM[45095] = 8'b11111011;
DRAM[45096] = 8'b11111101;
DRAM[45097] = 8'b11111110;
DRAM[45098] = 8'b11111110;
DRAM[45099] = 8'b11111111;
DRAM[45100] = 8'b11111111;
DRAM[45101] = 8'b11111110;
DRAM[45102] = 8'b11111110;
DRAM[45103] = 8'b11111101;
DRAM[45104] = 8'b11111111;
DRAM[45105] = 8'b11111110;
DRAM[45106] = 8'b11111101;
DRAM[45107] = 8'b11111101;
DRAM[45108] = 8'b11111101;
DRAM[45109] = 8'b11111101;
DRAM[45110] = 8'b11111010;
DRAM[45111] = 8'b11111000;
DRAM[45112] = 8'b11111000;
DRAM[45113] = 8'b11110101;
DRAM[45114] = 8'b11110000;
DRAM[45115] = 8'b11101101;
DRAM[45116] = 8'b11101011;
DRAM[45117] = 8'b11101010;
DRAM[45118] = 8'b11101000;
DRAM[45119] = 8'b11100110;
DRAM[45120] = 8'b11011100;
DRAM[45121] = 8'b11011001;
DRAM[45122] = 8'b11010010;
DRAM[45123] = 8'b11000111;
DRAM[45124] = 8'b10111100;
DRAM[45125] = 8'b10111000;
DRAM[45126] = 8'b10111011;
DRAM[45127] = 8'b10111111;
DRAM[45128] = 8'b10101000;
DRAM[45129] = 8'b10101011;
DRAM[45130] = 8'b10110101;
DRAM[45131] = 8'b10111110;
DRAM[45132] = 8'b10110110;
DRAM[45133] = 8'b10100100;
DRAM[45134] = 8'b10011101;
DRAM[45135] = 8'b10100010;
DRAM[45136] = 8'b10101010;
DRAM[45137] = 8'b10101000;
DRAM[45138] = 8'b10100110;
DRAM[45139] = 8'b10100000;
DRAM[45140] = 8'b10010111;
DRAM[45141] = 8'b10001110;
DRAM[45142] = 8'b10001010;
DRAM[45143] = 8'b10001011;
DRAM[45144] = 8'b10000110;
DRAM[45145] = 8'b10000011;
DRAM[45146] = 8'b10000001;
DRAM[45147] = 8'b10000011;
DRAM[45148] = 8'b10000111;
DRAM[45149] = 8'b10000111;
DRAM[45150] = 8'b10000011;
DRAM[45151] = 8'b1111111;
DRAM[45152] = 8'b10000101;
DRAM[45153] = 8'b10001011;
DRAM[45154] = 8'b10010011;
DRAM[45155] = 8'b10011011;
DRAM[45156] = 8'b10100011;
DRAM[45157] = 8'b10101001;
DRAM[45158] = 8'b10101010;
DRAM[45159] = 8'b10101000;
DRAM[45160] = 8'b10011010;
DRAM[45161] = 8'b10001011;
DRAM[45162] = 8'b1110110;
DRAM[45163] = 8'b1110000;
DRAM[45164] = 8'b10001001;
DRAM[45165] = 8'b10101111;
DRAM[45166] = 8'b11000101;
DRAM[45167] = 8'b11001000;
DRAM[45168] = 8'b10110110;
DRAM[45169] = 8'b10110000;
DRAM[45170] = 8'b10101100;
DRAM[45171] = 8'b10110010;
DRAM[45172] = 8'b11000000;
DRAM[45173] = 8'b11000101;
DRAM[45174] = 8'b10110111;
DRAM[45175] = 8'b10100100;
DRAM[45176] = 8'b10110011;
DRAM[45177] = 8'b10011000;
DRAM[45178] = 8'b10011010;
DRAM[45179] = 8'b10011011;
DRAM[45180] = 8'b10000001;
DRAM[45181] = 8'b1111111;
DRAM[45182] = 8'b10001000;
DRAM[45183] = 8'b1111001;
DRAM[45184] = 8'b1101101;
DRAM[45185] = 8'b1110011;
DRAM[45186] = 8'b1101011;
DRAM[45187] = 8'b1010111;
DRAM[45188] = 8'b1001111;
DRAM[45189] = 8'b1010010;
DRAM[45190] = 8'b1001100;
DRAM[45191] = 8'b111101;
DRAM[45192] = 8'b100100;
DRAM[45193] = 8'b11110;
DRAM[45194] = 8'b10110;
DRAM[45195] = 8'b10001;
DRAM[45196] = 8'b1110;
DRAM[45197] = 8'b1001;
DRAM[45198] = 8'b11;
DRAM[45199] = 8'b0;
DRAM[45200] = 8'b0;
DRAM[45201] = 8'b10;
DRAM[45202] = 8'b100;
DRAM[45203] = 8'b11;
DRAM[45204] = 8'b1;
DRAM[45205] = 8'b10;
DRAM[45206] = 8'b10;
DRAM[45207] = 8'b10;
DRAM[45208] = 8'b0;
DRAM[45209] = 8'b1;
DRAM[45210] = 8'b1;
DRAM[45211] = 8'b11;
DRAM[45212] = 8'b1101;
DRAM[45213] = 8'b11000;
DRAM[45214] = 8'b11101;
DRAM[45215] = 8'b11011;
DRAM[45216] = 8'b101010;
DRAM[45217] = 8'b101010;
DRAM[45218] = 8'b110101;
DRAM[45219] = 8'b1000111;
DRAM[45220] = 8'b1010010;
DRAM[45221] = 8'b1010110;
DRAM[45222] = 8'b1100010;
DRAM[45223] = 8'b1110001;
DRAM[45224] = 8'b1111110;
DRAM[45225] = 8'b10000000;
DRAM[45226] = 8'b10001011;
DRAM[45227] = 8'b10011011;
DRAM[45228] = 8'b10100000;
DRAM[45229] = 8'b10100010;
DRAM[45230] = 8'b10110100;
DRAM[45231] = 8'b11001100;
DRAM[45232] = 8'b11011101;
DRAM[45233] = 8'b11010110;
DRAM[45234] = 8'b11010010;
DRAM[45235] = 8'b11011011;
DRAM[45236] = 8'b11100110;
DRAM[45237] = 8'b11100001;
DRAM[45238] = 8'b11001010;
DRAM[45239] = 8'b10110010;
DRAM[45240] = 8'b11000001;
DRAM[45241] = 8'b11011011;
DRAM[45242] = 8'b11110011;
DRAM[45243] = 8'b11111001;
DRAM[45244] = 8'b11111001;
DRAM[45245] = 8'b11111011;
DRAM[45246] = 8'b11111000;
DRAM[45247] = 8'b11110001;
DRAM[45248] = 8'b11101001;
DRAM[45249] = 8'b11100100;
DRAM[45250] = 8'b11100000;
DRAM[45251] = 8'b11011100;
DRAM[45252] = 8'b11001111;
DRAM[45253] = 8'b10111101;
DRAM[45254] = 8'b10110011;
DRAM[45255] = 8'b10110010;
DRAM[45256] = 8'b10110001;
DRAM[45257] = 8'b10101101;
DRAM[45258] = 8'b10100101;
DRAM[45259] = 8'b10100011;
DRAM[45260] = 8'b10101101;
DRAM[45261] = 8'b10110101;
DRAM[45262] = 8'b10101000;
DRAM[45263] = 8'b10010011;
DRAM[45264] = 8'b10011100;
DRAM[45265] = 8'b10011001;
DRAM[45266] = 8'b10010101;
DRAM[45267] = 8'b10010010;
DRAM[45268] = 8'b10010001;
DRAM[45269] = 8'b10010001;
DRAM[45270] = 8'b10001111;
DRAM[45271] = 8'b10001110;
DRAM[45272] = 8'b10001011;
DRAM[45273] = 8'b10001001;
DRAM[45274] = 8'b10000111;
DRAM[45275] = 8'b10000110;
DRAM[45276] = 8'b10000111;
DRAM[45277] = 8'b10000111;
DRAM[45278] = 8'b10000110;
DRAM[45279] = 8'b10000101;
DRAM[45280] = 8'b10000010;
DRAM[45281] = 8'b10000001;
DRAM[45282] = 8'b10000000;
DRAM[45283] = 8'b10000000;
DRAM[45284] = 8'b1111111;
DRAM[45285] = 8'b1111110;
DRAM[45286] = 8'b1111101;
DRAM[45287] = 8'b1111101;
DRAM[45288] = 8'b1111100;
DRAM[45289] = 8'b1111100;
DRAM[45290] = 8'b1111101;
DRAM[45291] = 8'b1111101;
DRAM[45292] = 8'b1111111;
DRAM[45293] = 8'b10000001;
DRAM[45294] = 8'b10000010;
DRAM[45295] = 8'b10000011;
DRAM[45296] = 8'b10000110;
DRAM[45297] = 8'b10000110;
DRAM[45298] = 8'b10000111;
DRAM[45299] = 8'b10001000;
DRAM[45300] = 8'b10001000;
DRAM[45301] = 8'b10001000;
DRAM[45302] = 8'b10000111;
DRAM[45303] = 8'b10000111;
DRAM[45304] = 8'b10000111;
DRAM[45305] = 8'b10001000;
DRAM[45306] = 8'b10001010;
DRAM[45307] = 8'b10001011;
DRAM[45308] = 8'b10001100;
DRAM[45309] = 8'b10001011;
DRAM[45310] = 8'b10001011;
DRAM[45311] = 8'b10001010;
DRAM[45312] = 8'b10010001;
DRAM[45313] = 8'b10010000;
DRAM[45314] = 8'b10010000;
DRAM[45315] = 8'b10010000;
DRAM[45316] = 8'b10010000;
DRAM[45317] = 8'b10010001;
DRAM[45318] = 8'b10010010;
DRAM[45319] = 8'b10010011;
DRAM[45320] = 8'b10010011;
DRAM[45321] = 8'b10010100;
DRAM[45322] = 8'b10010101;
DRAM[45323] = 8'b10010110;
DRAM[45324] = 8'b10010111;
DRAM[45325] = 8'b10010111;
DRAM[45326] = 8'b10010111;
DRAM[45327] = 8'b10010111;
DRAM[45328] = 8'b10011000;
DRAM[45329] = 8'b10011000;
DRAM[45330] = 8'b10011001;
DRAM[45331] = 8'b10011001;
DRAM[45332] = 8'b10011010;
DRAM[45333] = 8'b10011011;
DRAM[45334] = 8'b10011100;
DRAM[45335] = 8'b10011100;
DRAM[45336] = 8'b10011110;
DRAM[45337] = 8'b10011100;
DRAM[45338] = 8'b10011011;
DRAM[45339] = 8'b10011101;
DRAM[45340] = 8'b10100000;
DRAM[45341] = 8'b10100001;
DRAM[45342] = 8'b10100000;
DRAM[45343] = 8'b10011110;
DRAM[45344] = 8'b10100011;
DRAM[45345] = 8'b10101001;
DRAM[45346] = 8'b10111110;
DRAM[45347] = 8'b11011100;
DRAM[45348] = 8'b11110100;
DRAM[45349] = 8'b11111110;
DRAM[45350] = 8'b11111111;
DRAM[45351] = 8'b11111111;
DRAM[45352] = 8'b11111101;
DRAM[45353] = 8'b11111110;
DRAM[45354] = 8'b11111110;
DRAM[45355] = 8'b11111111;
DRAM[45356] = 8'b11111111;
DRAM[45357] = 8'b11111110;
DRAM[45358] = 8'b11111110;
DRAM[45359] = 8'b11111101;
DRAM[45360] = 8'b11111011;
DRAM[45361] = 8'b11111010;
DRAM[45362] = 8'b11111001;
DRAM[45363] = 8'b11111001;
DRAM[45364] = 8'b11111001;
DRAM[45365] = 8'b11110111;
DRAM[45366] = 8'b11110100;
DRAM[45367] = 8'b11110001;
DRAM[45368] = 8'b11110000;
DRAM[45369] = 8'b11101110;
DRAM[45370] = 8'b11101100;
DRAM[45371] = 8'b11101011;
DRAM[45372] = 8'b11101001;
DRAM[45373] = 8'b11100110;
DRAM[45374] = 8'b11100010;
DRAM[45375] = 8'b11011110;
DRAM[45376] = 8'b11100110;
DRAM[45377] = 8'b11011011;
DRAM[45378] = 8'b11001101;
DRAM[45379] = 8'b11000101;
DRAM[45380] = 8'b11000010;
DRAM[45381] = 8'b10111011;
DRAM[45382] = 8'b10110000;
DRAM[45383] = 8'b10100110;
DRAM[45384] = 8'b10110000;
DRAM[45385] = 8'b10101101;
DRAM[45386] = 8'b10101111;
DRAM[45387] = 8'b10110011;
DRAM[45388] = 8'b10101110;
DRAM[45389] = 8'b10100101;
DRAM[45390] = 8'b10101000;
DRAM[45391] = 8'b10110011;
DRAM[45392] = 8'b10111010;
DRAM[45393] = 8'b10101100;
DRAM[45394] = 8'b10011110;
DRAM[45395] = 8'b10011100;
DRAM[45396] = 8'b10100000;
DRAM[45397] = 8'b10011110;
DRAM[45398] = 8'b10010010;
DRAM[45399] = 8'b10000111;
DRAM[45400] = 8'b10000111;
DRAM[45401] = 8'b10001001;
DRAM[45402] = 8'b10001011;
DRAM[45403] = 8'b10001010;
DRAM[45404] = 8'b10000110;
DRAM[45405] = 8'b10000011;
DRAM[45406] = 8'b10000010;
DRAM[45407] = 8'b10000010;
DRAM[45408] = 8'b10001100;
DRAM[45409] = 8'b10001101;
DRAM[45410] = 8'b10001111;
DRAM[45411] = 8'b10010100;
DRAM[45412] = 8'b10011100;
DRAM[45413] = 8'b10100111;
DRAM[45414] = 8'b10101111;
DRAM[45415] = 8'b10110010;
DRAM[45416] = 8'b10011101;
DRAM[45417] = 8'b10010010;
DRAM[45418] = 8'b1111111;
DRAM[45419] = 8'b1110001;
DRAM[45420] = 8'b1110101;
DRAM[45421] = 8'b10001011;
DRAM[45422] = 8'b10100101;
DRAM[45423] = 8'b10110100;
DRAM[45424] = 8'b11000000;
DRAM[45425] = 8'b11000010;
DRAM[45426] = 8'b11000001;
DRAM[45427] = 8'b10111110;
DRAM[45428] = 8'b10111101;
DRAM[45429] = 8'b10111101;
DRAM[45430] = 8'b10111000;
DRAM[45431] = 8'b10110001;
DRAM[45432] = 8'b10100011;
DRAM[45433] = 8'b10001110;
DRAM[45434] = 8'b10010010;
DRAM[45435] = 8'b10010011;
DRAM[45436] = 8'b10000001;
DRAM[45437] = 8'b10000111;
DRAM[45438] = 8'b10010000;
DRAM[45439] = 8'b1111111;
DRAM[45440] = 8'b1101111;
DRAM[45441] = 8'b1101101;
DRAM[45442] = 8'b1100000;
DRAM[45443] = 8'b1010011;
DRAM[45444] = 8'b1010011;
DRAM[45445] = 8'b1010101;
DRAM[45446] = 8'b1000011;
DRAM[45447] = 8'b101010;
DRAM[45448] = 8'b11010;
DRAM[45449] = 8'b10110;
DRAM[45450] = 8'b10010;
DRAM[45451] = 8'b1111;
DRAM[45452] = 8'b1101;
DRAM[45453] = 8'b1000;
DRAM[45454] = 8'b10;
DRAM[45455] = 8'b0;
DRAM[45456] = 8'b0;
DRAM[45457] = 8'b0;
DRAM[45458] = 8'b0;
DRAM[45459] = 8'b0;
DRAM[45460] = 8'b0;
DRAM[45461] = 8'b0;
DRAM[45462] = 8'b11;
DRAM[45463] = 8'b101;
DRAM[45464] = 8'b10;
DRAM[45465] = 8'b101;
DRAM[45466] = 8'b111;
DRAM[45467] = 8'b1001;
DRAM[45468] = 8'b10000;
DRAM[45469] = 8'b11001;
DRAM[45470] = 8'b11100;
DRAM[45471] = 8'b11010;
DRAM[45472] = 8'b100111;
DRAM[45473] = 8'b101011;
DRAM[45474] = 8'b111010;
DRAM[45475] = 8'b1001011;
DRAM[45476] = 8'b1010010;
DRAM[45477] = 8'b1010101;
DRAM[45478] = 8'b1100011;
DRAM[45479] = 8'b1110101;
DRAM[45480] = 8'b1111110;
DRAM[45481] = 8'b1111100;
DRAM[45482] = 8'b10000100;
DRAM[45483] = 8'b10010110;
DRAM[45484] = 8'b10100100;
DRAM[45485] = 8'b10101101;
DRAM[45486] = 8'b10111101;
DRAM[45487] = 8'b11010000;
DRAM[45488] = 8'b11100110;
DRAM[45489] = 8'b11100010;
DRAM[45490] = 8'b11011110;
DRAM[45491] = 8'b11011111;
DRAM[45492] = 8'b11100011;
DRAM[45493] = 8'b11011110;
DRAM[45494] = 8'b11001001;
DRAM[45495] = 8'b10110010;
DRAM[45496] = 8'b11000101;
DRAM[45497] = 8'b11011110;
DRAM[45498] = 8'b11110100;
DRAM[45499] = 8'b11111010;
DRAM[45500] = 8'b11111010;
DRAM[45501] = 8'b11111100;
DRAM[45502] = 8'b11111001;
DRAM[45503] = 8'b11110011;
DRAM[45504] = 8'b11101111;
DRAM[45505] = 8'b11101001;
DRAM[45506] = 8'b11100100;
DRAM[45507] = 8'b11100000;
DRAM[45508] = 8'b11010100;
DRAM[45509] = 8'b11000010;
DRAM[45510] = 8'b10110101;
DRAM[45511] = 8'b10110010;
DRAM[45512] = 8'b10101111;
DRAM[45513] = 8'b10101100;
DRAM[45514] = 8'b10100110;
DRAM[45515] = 8'b10100100;
DRAM[45516] = 8'b10101000;
DRAM[45517] = 8'b10101011;
DRAM[45518] = 8'b10100101;
DRAM[45519] = 8'b10011100;
DRAM[45520] = 8'b10011001;
DRAM[45521] = 8'b10010110;
DRAM[45522] = 8'b10010010;
DRAM[45523] = 8'b10010000;
DRAM[45524] = 8'b10001111;
DRAM[45525] = 8'b10001110;
DRAM[45526] = 8'b10001100;
DRAM[45527] = 8'b10001010;
DRAM[45528] = 8'b10001001;
DRAM[45529] = 8'b10000111;
DRAM[45530] = 8'b10000101;
DRAM[45531] = 8'b10000100;
DRAM[45532] = 8'b10000101;
DRAM[45533] = 8'b10000101;
DRAM[45534] = 8'b10000100;
DRAM[45535] = 8'b10000011;
DRAM[45536] = 8'b10000001;
DRAM[45537] = 8'b10000001;
DRAM[45538] = 8'b10000000;
DRAM[45539] = 8'b1111111;
DRAM[45540] = 8'b1111110;
DRAM[45541] = 8'b1111101;
DRAM[45542] = 8'b1111101;
DRAM[45543] = 8'b1111100;
DRAM[45544] = 8'b1111101;
DRAM[45545] = 8'b1111101;
DRAM[45546] = 8'b1111101;
DRAM[45547] = 8'b1111110;
DRAM[45548] = 8'b1111111;
DRAM[45549] = 8'b10000001;
DRAM[45550] = 8'b10000010;
DRAM[45551] = 8'b10000011;
DRAM[45552] = 8'b10000110;
DRAM[45553] = 8'b10000110;
DRAM[45554] = 8'b10000111;
DRAM[45555] = 8'b10000111;
DRAM[45556] = 8'b10001000;
DRAM[45557] = 8'b10001000;
DRAM[45558] = 8'b10001000;
DRAM[45559] = 8'b10000111;
DRAM[45560] = 8'b10001000;
DRAM[45561] = 8'b10001001;
DRAM[45562] = 8'b10001010;
DRAM[45563] = 8'b10001011;
DRAM[45564] = 8'b10001100;
DRAM[45565] = 8'b10001011;
DRAM[45566] = 8'b10001011;
DRAM[45567] = 8'b10001010;
DRAM[45568] = 8'b10010000;
DRAM[45569] = 8'b10010000;
DRAM[45570] = 8'b10010000;
DRAM[45571] = 8'b10010000;
DRAM[45572] = 8'b10010000;
DRAM[45573] = 8'b10010001;
DRAM[45574] = 8'b10010010;
DRAM[45575] = 8'b10010010;
DRAM[45576] = 8'b10010100;
DRAM[45577] = 8'b10010100;
DRAM[45578] = 8'b10010101;
DRAM[45579] = 8'b10010110;
DRAM[45580] = 8'b10010110;
DRAM[45581] = 8'b10010110;
DRAM[45582] = 8'b10010101;
DRAM[45583] = 8'b10010101;
DRAM[45584] = 8'b10010111;
DRAM[45585] = 8'b10010111;
DRAM[45586] = 8'b10011000;
DRAM[45587] = 8'b10011001;
DRAM[45588] = 8'b10011010;
DRAM[45589] = 8'b10011010;
DRAM[45590] = 8'b10011011;
DRAM[45591] = 8'b10011011;
DRAM[45592] = 8'b10011100;
DRAM[45593] = 8'b10011011;
DRAM[45594] = 8'b10011010;
DRAM[45595] = 8'b10011011;
DRAM[45596] = 8'b10011101;
DRAM[45597] = 8'b10011111;
DRAM[45598] = 8'b10100000;
DRAM[45599] = 8'b10011111;
DRAM[45600] = 8'b10100110;
DRAM[45601] = 8'b10110011;
DRAM[45602] = 8'b11001011;
DRAM[45603] = 8'b11100111;
DRAM[45604] = 8'b11111001;
DRAM[45605] = 8'b11111111;
DRAM[45606] = 8'b11111111;
DRAM[45607] = 8'b11111111;
DRAM[45608] = 8'b11111101;
DRAM[45609] = 8'b11111110;
DRAM[45610] = 8'b11111110;
DRAM[45611] = 8'b11111111;
DRAM[45612] = 8'b11111111;
DRAM[45613] = 8'b11111110;
DRAM[45614] = 8'b11111110;
DRAM[45615] = 8'b11111101;
DRAM[45616] = 8'b11111100;
DRAM[45617] = 8'b11111011;
DRAM[45618] = 8'b11111011;
DRAM[45619] = 8'b11111011;
DRAM[45620] = 8'b11111011;
DRAM[45621] = 8'b11111000;
DRAM[45622] = 8'b11110100;
DRAM[45623] = 8'b11110000;
DRAM[45624] = 8'b11101100;
DRAM[45625] = 8'b11101011;
DRAM[45626] = 8'b11101010;
DRAM[45627] = 8'b11101000;
DRAM[45628] = 8'b11100101;
DRAM[45629] = 8'b11011111;
DRAM[45630] = 8'b11011000;
DRAM[45631] = 8'b11010011;
DRAM[45632] = 8'b11000111;
DRAM[45633] = 8'b11000011;
DRAM[45634] = 8'b11000010;
DRAM[45635] = 8'b11000111;
DRAM[45636] = 8'b11001111;
DRAM[45637] = 8'b11010000;
DRAM[45638] = 8'b11001000;
DRAM[45639] = 8'b10111111;
DRAM[45640] = 8'b11000100;
DRAM[45641] = 8'b10111100;
DRAM[45642] = 8'b10110110;
DRAM[45643] = 8'b10110010;
DRAM[45644] = 8'b10101001;
DRAM[45645] = 8'b10100000;
DRAM[45646] = 8'b10100011;
DRAM[45647] = 8'b10101100;
DRAM[45648] = 8'b10110010;
DRAM[45649] = 8'b10110000;
DRAM[45650] = 8'b10101100;
DRAM[45651] = 8'b10100110;
DRAM[45652] = 8'b10100000;
DRAM[45653] = 8'b10011101;
DRAM[45654] = 8'b10011010;
DRAM[45655] = 8'b10011001;
DRAM[45656] = 8'b10000111;
DRAM[45657] = 8'b10001100;
DRAM[45658] = 8'b10001111;
DRAM[45659] = 8'b10001010;
DRAM[45660] = 8'b10000001;
DRAM[45661] = 8'b1111011;
DRAM[45662] = 8'b1111110;
DRAM[45663] = 8'b10000011;
DRAM[45664] = 8'b10010111;
DRAM[45665] = 8'b10010010;
DRAM[45666] = 8'b10001100;
DRAM[45667] = 8'b10001010;
DRAM[45668] = 8'b10001111;
DRAM[45669] = 8'b10011010;
DRAM[45670] = 8'b10100111;
DRAM[45671] = 8'b10110001;
DRAM[45672] = 8'b10100010;
DRAM[45673] = 8'b10011101;
DRAM[45674] = 8'b10001011;
DRAM[45675] = 8'b1101100;
DRAM[45676] = 8'b1010011;
DRAM[45677] = 8'b1011110;
DRAM[45678] = 8'b10010000;
DRAM[45679] = 8'b11000001;
DRAM[45680] = 8'b11000001;
DRAM[45681] = 8'b11000100;
DRAM[45682] = 8'b11000010;
DRAM[45683] = 8'b10111100;
DRAM[45684] = 8'b10110111;
DRAM[45685] = 8'b10110101;
DRAM[45686] = 8'b10110011;
DRAM[45687] = 8'b10101111;
DRAM[45688] = 8'b10011111;
DRAM[45689] = 8'b10010010;
DRAM[45690] = 8'b10010011;
DRAM[45691] = 8'b10001110;
DRAM[45692] = 8'b10000001;
DRAM[45693] = 8'b10001011;
DRAM[45694] = 8'b10010000;
DRAM[45695] = 8'b1111010;
DRAM[45696] = 8'b1101110;
DRAM[45697] = 8'b1101101;
DRAM[45698] = 8'b1100010;
DRAM[45699] = 8'b1010101;
DRAM[45700] = 8'b1010010;
DRAM[45701] = 8'b1010000;
DRAM[45702] = 8'b111101;
DRAM[45703] = 8'b100101;
DRAM[45704] = 8'b11010;
DRAM[45705] = 8'b11001;
DRAM[45706] = 8'b11000;
DRAM[45707] = 8'b10110;
DRAM[45708] = 8'b10010;
DRAM[45709] = 8'b1110;
DRAM[45710] = 8'b1010;
DRAM[45711] = 8'b111;
DRAM[45712] = 8'b100;
DRAM[45713] = 8'b11;
DRAM[45714] = 8'b1;
DRAM[45715] = 8'b0;
DRAM[45716] = 8'b0;
DRAM[45717] = 8'b10;
DRAM[45718] = 8'b1001;
DRAM[45719] = 8'b1110;
DRAM[45720] = 8'b1001;
DRAM[45721] = 8'b1111;
DRAM[45722] = 8'b10011;
DRAM[45723] = 8'b10011;
DRAM[45724] = 8'b10101;
DRAM[45725] = 8'b11010;
DRAM[45726] = 8'b11100;
DRAM[45727] = 8'b11011;
DRAM[45728] = 8'b11100;
DRAM[45729] = 8'b100100;
DRAM[45730] = 8'b110101;
DRAM[45731] = 8'b1000100;
DRAM[45732] = 8'b1001001;
DRAM[45733] = 8'b1001100;
DRAM[45734] = 8'b1011011;
DRAM[45735] = 8'b1101110;
DRAM[45736] = 8'b1111001;
DRAM[45737] = 8'b1110011;
DRAM[45738] = 8'b1111000;
DRAM[45739] = 8'b10001011;
DRAM[45740] = 8'b10100001;
DRAM[45741] = 8'b10110010;
DRAM[45742] = 8'b11000001;
DRAM[45743] = 8'b11001101;
DRAM[45744] = 8'b11011001;
DRAM[45745] = 8'b11011001;
DRAM[45746] = 8'b11011011;
DRAM[45747] = 8'b11011111;
DRAM[45748] = 8'b11100001;
DRAM[45749] = 8'b11011101;
DRAM[45750] = 8'b11010001;
DRAM[45751] = 8'b11000101;
DRAM[45752] = 8'b11001110;
DRAM[45753] = 8'b11100011;
DRAM[45754] = 8'b11110110;
DRAM[45755] = 8'b11111011;
DRAM[45756] = 8'b11111011;
DRAM[45757] = 8'b11111101;
DRAM[45758] = 8'b11111011;
DRAM[45759] = 8'b11110110;
DRAM[45760] = 8'b11110010;
DRAM[45761] = 8'b11101100;
DRAM[45762] = 8'b11100101;
DRAM[45763] = 8'b11100000;
DRAM[45764] = 8'b11010110;
DRAM[45765] = 8'b11000110;
DRAM[45766] = 8'b10110110;
DRAM[45767] = 8'b10101101;
DRAM[45768] = 8'b10101101;
DRAM[45769] = 8'b10101001;
DRAM[45770] = 8'b10100110;
DRAM[45771] = 8'b10100101;
DRAM[45772] = 8'b10100010;
DRAM[45773] = 8'b10011111;
DRAM[45774] = 8'b10100000;
DRAM[45775] = 8'b10100100;
DRAM[45776] = 8'b10010101;
DRAM[45777] = 8'b10010011;
DRAM[45778] = 8'b10010000;
DRAM[45779] = 8'b10001110;
DRAM[45780] = 8'b10001101;
DRAM[45781] = 8'b10001011;
DRAM[45782] = 8'b10001000;
DRAM[45783] = 8'b10000110;
DRAM[45784] = 8'b10000111;
DRAM[45785] = 8'b10000101;
DRAM[45786] = 8'b10000011;
DRAM[45787] = 8'b10000010;
DRAM[45788] = 8'b10000011;
DRAM[45789] = 8'b10000011;
DRAM[45790] = 8'b10000010;
DRAM[45791] = 8'b10000001;
DRAM[45792] = 8'b10000000;
DRAM[45793] = 8'b10000000;
DRAM[45794] = 8'b1111111;
DRAM[45795] = 8'b1111111;
DRAM[45796] = 8'b1111110;
DRAM[45797] = 8'b1111101;
DRAM[45798] = 8'b1111101;
DRAM[45799] = 8'b1111100;
DRAM[45800] = 8'b1111101;
DRAM[45801] = 8'b1111101;
DRAM[45802] = 8'b1111101;
DRAM[45803] = 8'b1111110;
DRAM[45804] = 8'b1111111;
DRAM[45805] = 8'b10000001;
DRAM[45806] = 8'b10000010;
DRAM[45807] = 8'b10000011;
DRAM[45808] = 8'b10000110;
DRAM[45809] = 8'b10000110;
DRAM[45810] = 8'b10000110;
DRAM[45811] = 8'b10000111;
DRAM[45812] = 8'b10000111;
DRAM[45813] = 8'b10001000;
DRAM[45814] = 8'b10001000;
DRAM[45815] = 8'b10001000;
DRAM[45816] = 8'b10001001;
DRAM[45817] = 8'b10001001;
DRAM[45818] = 8'b10001010;
DRAM[45819] = 8'b10001011;
DRAM[45820] = 8'b10001011;
DRAM[45821] = 8'b10001011;
DRAM[45822] = 8'b10001011;
DRAM[45823] = 8'b10001010;
DRAM[45824] = 8'b10010000;
DRAM[45825] = 8'b10010000;
DRAM[45826] = 8'b10001111;
DRAM[45827] = 8'b10001111;
DRAM[45828] = 8'b10010000;
DRAM[45829] = 8'b10010000;
DRAM[45830] = 8'b10010001;
DRAM[45831] = 8'b10010010;
DRAM[45832] = 8'b10010101;
DRAM[45833] = 8'b10010101;
DRAM[45834] = 8'b10010110;
DRAM[45835] = 8'b10010110;
DRAM[45836] = 8'b10010110;
DRAM[45837] = 8'b10010101;
DRAM[45838] = 8'b10010100;
DRAM[45839] = 8'b10010100;
DRAM[45840] = 8'b10010110;
DRAM[45841] = 8'b10010111;
DRAM[45842] = 8'b10010111;
DRAM[45843] = 8'b10011000;
DRAM[45844] = 8'b10011001;
DRAM[45845] = 8'b10011010;
DRAM[45846] = 8'b10011010;
DRAM[45847] = 8'b10011010;
DRAM[45848] = 8'b10011010;
DRAM[45849] = 8'b10011001;
DRAM[45850] = 8'b10011001;
DRAM[45851] = 8'b10011001;
DRAM[45852] = 8'b10011100;
DRAM[45853] = 8'b10011110;
DRAM[45854] = 8'b10100001;
DRAM[45855] = 8'b10100010;
DRAM[45856] = 8'b10101110;
DRAM[45857] = 8'b10111111;
DRAM[45858] = 8'b11011001;
DRAM[45859] = 8'b11101111;
DRAM[45860] = 8'b11111011;
DRAM[45861] = 8'b11111110;
DRAM[45862] = 8'b11111110;
DRAM[45863] = 8'b11111111;
DRAM[45864] = 8'b11111101;
DRAM[45865] = 8'b11111110;
DRAM[45866] = 8'b11111110;
DRAM[45867] = 8'b11111111;
DRAM[45868] = 8'b11111111;
DRAM[45869] = 8'b11111110;
DRAM[45870] = 8'b11111110;
DRAM[45871] = 8'b11111101;
DRAM[45872] = 8'b11111110;
DRAM[45873] = 8'b11111101;
DRAM[45874] = 8'b11111101;
DRAM[45875] = 8'b11111101;
DRAM[45876] = 8'b11111100;
DRAM[45877] = 8'b11111001;
DRAM[45878] = 8'b11110100;
DRAM[45879] = 8'b11110000;
DRAM[45880] = 8'b11110000;
DRAM[45881] = 8'b11101110;
DRAM[45882] = 8'b11101010;
DRAM[45883] = 8'b11100110;
DRAM[45884] = 8'b11100010;
DRAM[45885] = 8'b11011100;
DRAM[45886] = 8'b11010100;
DRAM[45887] = 8'b11001111;
DRAM[45888] = 8'b11001100;
DRAM[45889] = 8'b11010010;
DRAM[45890] = 8'b11011000;
DRAM[45891] = 8'b11011000;
DRAM[45892] = 8'b11010010;
DRAM[45893] = 8'b11001100;
DRAM[45894] = 8'b11001001;
DRAM[45895] = 8'b11001001;
DRAM[45896] = 8'b11001010;
DRAM[45897] = 8'b11000100;
DRAM[45898] = 8'b10111110;
DRAM[45899] = 8'b10111000;
DRAM[45900] = 8'b10101101;
DRAM[45901] = 8'b10100000;
DRAM[45902] = 8'b10011010;
DRAM[45903] = 8'b10011011;
DRAM[45904] = 8'b10100101;
DRAM[45905] = 8'b10101111;
DRAM[45906] = 8'b10110101;
DRAM[45907] = 8'b10101111;
DRAM[45908] = 8'b10100110;
DRAM[45909] = 8'b10100000;
DRAM[45910] = 8'b10011111;
DRAM[45911] = 8'b10100000;
DRAM[45912] = 8'b10001101;
DRAM[45913] = 8'b10001111;
DRAM[45914] = 8'b10001111;
DRAM[45915] = 8'b10001000;
DRAM[45916] = 8'b1111111;
DRAM[45917] = 8'b1111100;
DRAM[45918] = 8'b10000001;
DRAM[45919] = 8'b10001000;
DRAM[45920] = 8'b10001111;
DRAM[45921] = 8'b10001001;
DRAM[45922] = 8'b10000011;
DRAM[45923] = 8'b10000010;
DRAM[45924] = 8'b10000110;
DRAM[45925] = 8'b10010000;
DRAM[45926] = 8'b10011111;
DRAM[45927] = 8'b10101100;
DRAM[45928] = 8'b10101001;
DRAM[45929] = 8'b10011011;
DRAM[45930] = 8'b10000110;
DRAM[45931] = 8'b1101111;
DRAM[45932] = 8'b1011101;
DRAM[45933] = 8'b1100101;
DRAM[45934] = 8'b10001101;
DRAM[45935] = 8'b10111000;
DRAM[45936] = 8'b10111100;
DRAM[45937] = 8'b10111000;
DRAM[45938] = 8'b10110011;
DRAM[45939] = 8'b10110001;
DRAM[45940] = 8'b10110101;
DRAM[45941] = 8'b10110111;
DRAM[45942] = 8'b10101110;
DRAM[45943] = 8'b10100001;
DRAM[45944] = 8'b10100000;
DRAM[45945] = 8'b10011010;
DRAM[45946] = 8'b10010111;
DRAM[45947] = 8'b10001101;
DRAM[45948] = 8'b10000100;
DRAM[45949] = 8'b10001110;
DRAM[45950] = 8'b10001110;
DRAM[45951] = 8'b1110110;
DRAM[45952] = 8'b1101010;
DRAM[45953] = 8'b1110000;
DRAM[45954] = 8'b1101011;
DRAM[45955] = 8'b1011001;
DRAM[45956] = 8'b1001011;
DRAM[45957] = 8'b1000101;
DRAM[45958] = 8'b111110;
DRAM[45959] = 8'b110100;
DRAM[45960] = 8'b100011;
DRAM[45961] = 8'b100010;
DRAM[45962] = 8'b11110;
DRAM[45963] = 8'b11010;
DRAM[45964] = 8'b10101;
DRAM[45965] = 8'b10010;
DRAM[45966] = 8'b10000;
DRAM[45967] = 8'b1111;
DRAM[45968] = 8'b1001;
DRAM[45969] = 8'b110;
DRAM[45970] = 8'b100;
DRAM[45971] = 8'b100;
DRAM[45972] = 8'b100;
DRAM[45973] = 8'b101;
DRAM[45974] = 8'b1011;
DRAM[45975] = 8'b10010;
DRAM[45976] = 8'b10001;
DRAM[45977] = 8'b10111;
DRAM[45978] = 8'b11010;
DRAM[45979] = 8'b10110;
DRAM[45980] = 8'b10100;
DRAM[45981] = 8'b10110;
DRAM[45982] = 8'b11001;
DRAM[45983] = 8'b11010;
DRAM[45984] = 8'b11000;
DRAM[45985] = 8'b11111;
DRAM[45986] = 8'b101101;
DRAM[45987] = 8'b111011;
DRAM[45988] = 8'b1000010;
DRAM[45989] = 8'b1001000;
DRAM[45990] = 8'b1010101;
DRAM[45991] = 8'b1100011;
DRAM[45992] = 8'b1110110;
DRAM[45993] = 8'b1110011;
DRAM[45994] = 8'b1110111;
DRAM[45995] = 8'b10000111;
DRAM[45996] = 8'b10011101;
DRAM[45997] = 8'b10110001;
DRAM[45998] = 8'b11000001;
DRAM[45999] = 8'b11001010;
DRAM[46000] = 8'b11000110;
DRAM[46001] = 8'b11000101;
DRAM[46002] = 8'b11001111;
DRAM[46003] = 8'b11011110;
DRAM[46004] = 8'b11011110;
DRAM[46005] = 8'b11010011;
DRAM[46006] = 8'b11001111;
DRAM[46007] = 8'b11010110;
DRAM[46008] = 8'b11011000;
DRAM[46009] = 8'b11101001;
DRAM[46010] = 8'b11111000;
DRAM[46011] = 8'b11111101;
DRAM[46012] = 8'b11111100;
DRAM[46013] = 8'b11111101;
DRAM[46014] = 8'b11111101;
DRAM[46015] = 8'b11111010;
DRAM[46016] = 8'b11110111;
DRAM[46017] = 8'b11110000;
DRAM[46018] = 8'b11101001;
DRAM[46019] = 8'b11100100;
DRAM[46020] = 8'b11011100;
DRAM[46021] = 8'b11001110;
DRAM[46022] = 8'b10111101;
DRAM[46023] = 8'b10110001;
DRAM[46024] = 8'b10101100;
DRAM[46025] = 8'b10100110;
DRAM[46026] = 8'b10100011;
DRAM[46027] = 8'b10100110;
DRAM[46028] = 8'b10100010;
DRAM[46029] = 8'b10011010;
DRAM[46030] = 8'b10011011;
DRAM[46031] = 8'b10100011;
DRAM[46032] = 8'b10010100;
DRAM[46033] = 8'b10010001;
DRAM[46034] = 8'b10001111;
DRAM[46035] = 8'b10001101;
DRAM[46036] = 8'b10001100;
DRAM[46037] = 8'b10001010;
DRAM[46038] = 8'b10000110;
DRAM[46039] = 8'b10000011;
DRAM[46040] = 8'b10000110;
DRAM[46041] = 8'b10000100;
DRAM[46042] = 8'b10000010;
DRAM[46043] = 8'b10000001;
DRAM[46044] = 8'b10000010;
DRAM[46045] = 8'b10000010;
DRAM[46046] = 8'b10000001;
DRAM[46047] = 8'b10000000;
DRAM[46048] = 8'b1111111;
DRAM[46049] = 8'b1111111;
DRAM[46050] = 8'b1111110;
DRAM[46051] = 8'b1111110;
DRAM[46052] = 8'b1111101;
DRAM[46053] = 8'b1111101;
DRAM[46054] = 8'b1111100;
DRAM[46055] = 8'b1111100;
DRAM[46056] = 8'b1111110;
DRAM[46057] = 8'b1111110;
DRAM[46058] = 8'b1111110;
DRAM[46059] = 8'b1111110;
DRAM[46060] = 8'b1111111;
DRAM[46061] = 8'b10000001;
DRAM[46062] = 8'b10000010;
DRAM[46063] = 8'b10000011;
DRAM[46064] = 8'b10000110;
DRAM[46065] = 8'b10000110;
DRAM[46066] = 8'b10000110;
DRAM[46067] = 8'b10000110;
DRAM[46068] = 8'b10000111;
DRAM[46069] = 8'b10001000;
DRAM[46070] = 8'b10001001;
DRAM[46071] = 8'b10001001;
DRAM[46072] = 8'b10001010;
DRAM[46073] = 8'b10001010;
DRAM[46074] = 8'b10001011;
DRAM[46075] = 8'b10001011;
DRAM[46076] = 8'b10001011;
DRAM[46077] = 8'b10001011;
DRAM[46078] = 8'b10001011;
DRAM[46079] = 8'b10001011;
DRAM[46080] = 8'b10010000;
DRAM[46081] = 8'b10001111;
DRAM[46082] = 8'b10001111;
DRAM[46083] = 8'b10001111;
DRAM[46084] = 8'b10001111;
DRAM[46085] = 8'b10010000;
DRAM[46086] = 8'b10010001;
DRAM[46087] = 8'b10010010;
DRAM[46088] = 8'b10010101;
DRAM[46089] = 8'b10010101;
DRAM[46090] = 8'b10010110;
DRAM[46091] = 8'b10010110;
DRAM[46092] = 8'b10010110;
DRAM[46093] = 8'b10010101;
DRAM[46094] = 8'b10010100;
DRAM[46095] = 8'b10010100;
DRAM[46096] = 8'b10010110;
DRAM[46097] = 8'b10010110;
DRAM[46098] = 8'b10010110;
DRAM[46099] = 8'b10010111;
DRAM[46100] = 8'b10011000;
DRAM[46101] = 8'b10011001;
DRAM[46102] = 8'b10011001;
DRAM[46103] = 8'b10011010;
DRAM[46104] = 8'b10011001;
DRAM[46105] = 8'b10011000;
DRAM[46106] = 8'b10011000;
DRAM[46107] = 8'b10011001;
DRAM[46108] = 8'b10011011;
DRAM[46109] = 8'b10011111;
DRAM[46110] = 8'b10100100;
DRAM[46111] = 8'b10101000;
DRAM[46112] = 8'b10111011;
DRAM[46113] = 8'b11001110;
DRAM[46114] = 8'b11100111;
DRAM[46115] = 8'b11110110;
DRAM[46116] = 8'b11111100;
DRAM[46117] = 8'b11111101;
DRAM[46118] = 8'b11111101;
DRAM[46119] = 8'b11111101;
DRAM[46120] = 8'b11111101;
DRAM[46121] = 8'b11111110;
DRAM[46122] = 8'b11111110;
DRAM[46123] = 8'b11111111;
DRAM[46124] = 8'b11111111;
DRAM[46125] = 8'b11111110;
DRAM[46126] = 8'b11111110;
DRAM[46127] = 8'b11111101;
DRAM[46128] = 8'b11111011;
DRAM[46129] = 8'b11111010;
DRAM[46130] = 8'b11111001;
DRAM[46131] = 8'b11111001;
DRAM[46132] = 8'b11111000;
DRAM[46133] = 8'b11110110;
DRAM[46134] = 8'b11110001;
DRAM[46135] = 8'b11101101;
DRAM[46136] = 8'b11110010;
DRAM[46137] = 8'b11101111;
DRAM[46138] = 8'b11101010;
DRAM[46139] = 8'b11100110;
DRAM[46140] = 8'b11100011;
DRAM[46141] = 8'b11100000;
DRAM[46142] = 8'b11011100;
DRAM[46143] = 8'b11011001;
DRAM[46144] = 8'b11100000;
DRAM[46145] = 8'b11100100;
DRAM[46146] = 8'b11100101;
DRAM[46147] = 8'b11011111;
DRAM[46148] = 8'b11010101;
DRAM[46149] = 8'b11001100;
DRAM[46150] = 8'b11001000;
DRAM[46151] = 8'b11001000;
DRAM[46152] = 8'b11000000;
DRAM[46153] = 8'b10111100;
DRAM[46154] = 8'b10111001;
DRAM[46155] = 8'b10111000;
DRAM[46156] = 8'b10110010;
DRAM[46157] = 8'b10101001;
DRAM[46158] = 8'b10100001;
DRAM[46159] = 8'b10011110;
DRAM[46160] = 8'b10101001;
DRAM[46161] = 8'b10101011;
DRAM[46162] = 8'b10101100;
DRAM[46163] = 8'b10101101;
DRAM[46164] = 8'b10110001;
DRAM[46165] = 8'b10101111;
DRAM[46166] = 8'b10100000;
DRAM[46167] = 8'b10001111;
DRAM[46168] = 8'b10010110;
DRAM[46169] = 8'b10010010;
DRAM[46170] = 8'b10001011;
DRAM[46171] = 8'b10000101;
DRAM[46172] = 8'b10000011;
DRAM[46173] = 8'b10000110;
DRAM[46174] = 8'b10001010;
DRAM[46175] = 8'b10001110;
DRAM[46176] = 8'b1111101;
DRAM[46177] = 8'b1111010;
DRAM[46178] = 8'b1111011;
DRAM[46179] = 8'b10000010;
DRAM[46180] = 8'b10000111;
DRAM[46181] = 8'b10001110;
DRAM[46182] = 8'b10011011;
DRAM[46183] = 8'b10101000;
DRAM[46184] = 8'b10101011;
DRAM[46185] = 8'b10010100;
DRAM[46186] = 8'b10000010;
DRAM[46187] = 8'b10000011;
DRAM[46188] = 8'b10001001;
DRAM[46189] = 8'b10000111;
DRAM[46190] = 8'b10000001;
DRAM[46191] = 8'b1111111;
DRAM[46192] = 8'b10110000;
DRAM[46193] = 8'b10110011;
DRAM[46194] = 8'b10110101;
DRAM[46195] = 8'b10110110;
DRAM[46196] = 8'b10111001;
DRAM[46197] = 8'b10110111;
DRAM[46198] = 8'b10101101;
DRAM[46199] = 8'b10100010;
DRAM[46200] = 8'b10011010;
DRAM[46201] = 8'b10011011;
DRAM[46202] = 8'b10010110;
DRAM[46203] = 8'b10001011;
DRAM[46204] = 8'b10000111;
DRAM[46205] = 8'b10001110;
DRAM[46206] = 8'b10001011;
DRAM[46207] = 8'b1111000;
DRAM[46208] = 8'b1101100;
DRAM[46209] = 8'b1101100;
DRAM[46210] = 8'b1100010;
DRAM[46211] = 8'b1010000;
DRAM[46212] = 8'b1000100;
DRAM[46213] = 8'b1000010;
DRAM[46214] = 8'b1000001;
DRAM[46215] = 8'b111100;
DRAM[46216] = 8'b101011;
DRAM[46217] = 8'b100101;
DRAM[46218] = 8'b11100;
DRAM[46219] = 8'b10100;
DRAM[46220] = 8'b10000;
DRAM[46221] = 8'b1110;
DRAM[46222] = 8'b1111;
DRAM[46223] = 8'b1111;
DRAM[46224] = 8'b1110;
DRAM[46225] = 8'b1010;
DRAM[46226] = 8'b1000;
DRAM[46227] = 8'b1010;
DRAM[46228] = 8'b1000;
DRAM[46229] = 8'b110;
DRAM[46230] = 8'b1001;
DRAM[46231] = 8'b10001;
DRAM[46232] = 8'b11000;
DRAM[46233] = 8'b11101;
DRAM[46234] = 8'b11101;
DRAM[46235] = 8'b11000;
DRAM[46236] = 8'b10100;
DRAM[46237] = 8'b10111;
DRAM[46238] = 8'b11010;
DRAM[46239] = 8'b11010;
DRAM[46240] = 8'b100011;
DRAM[46241] = 8'b100101;
DRAM[46242] = 8'b101101;
DRAM[46243] = 8'b111010;
DRAM[46244] = 8'b1000101;
DRAM[46245] = 8'b1001110;
DRAM[46246] = 8'b1010111;
DRAM[46247] = 8'b1011110;
DRAM[46248] = 8'b1110110;
DRAM[46249] = 8'b1111100;
DRAM[46250] = 8'b10000011;
DRAM[46251] = 8'b10001101;
DRAM[46252] = 8'b10011101;
DRAM[46253] = 8'b10110000;
DRAM[46254] = 8'b11000000;
DRAM[46255] = 8'b11001000;
DRAM[46256] = 8'b11000110;
DRAM[46257] = 8'b11000000;
DRAM[46258] = 8'b11001100;
DRAM[46259] = 8'b11100000;
DRAM[46260] = 8'b11011010;
DRAM[46261] = 8'b11000011;
DRAM[46262] = 8'b11000011;
DRAM[46263] = 8'b11011000;
DRAM[46264] = 8'b11100011;
DRAM[46265] = 8'b11101110;
DRAM[46266] = 8'b11111001;
DRAM[46267] = 8'b11111101;
DRAM[46268] = 8'b11111101;
DRAM[46269] = 8'b11111101;
DRAM[46270] = 8'b11111110;
DRAM[46271] = 8'b11111101;
DRAM[46272] = 8'b11111110;
DRAM[46273] = 8'b11111001;
DRAM[46274] = 8'b11110010;
DRAM[46275] = 8'b11101100;
DRAM[46276] = 8'b11100101;
DRAM[46277] = 8'b11011010;
DRAM[46278] = 8'b11001010;
DRAM[46279] = 8'b10111101;
DRAM[46280] = 8'b10101101;
DRAM[46281] = 8'b10100100;
DRAM[46282] = 8'b10100001;
DRAM[46283] = 8'b10100101;
DRAM[46284] = 8'b10100100;
DRAM[46285] = 8'b10011011;
DRAM[46286] = 8'b10011000;
DRAM[46287] = 8'b10011011;
DRAM[46288] = 8'b10010101;
DRAM[46289] = 8'b10010010;
DRAM[46290] = 8'b10001111;
DRAM[46291] = 8'b10001100;
DRAM[46292] = 8'b10001011;
DRAM[46293] = 8'b10001001;
DRAM[46294] = 8'b10000110;
DRAM[46295] = 8'b10000011;
DRAM[46296] = 8'b10000110;
DRAM[46297] = 8'b10000100;
DRAM[46298] = 8'b10000001;
DRAM[46299] = 8'b10000001;
DRAM[46300] = 8'b10000001;
DRAM[46301] = 8'b10000010;
DRAM[46302] = 8'b10000001;
DRAM[46303] = 8'b1111111;
DRAM[46304] = 8'b1111101;
DRAM[46305] = 8'b1111101;
DRAM[46306] = 8'b1111101;
DRAM[46307] = 8'b1111101;
DRAM[46308] = 8'b1111100;
DRAM[46309] = 8'b1111100;
DRAM[46310] = 8'b1111100;
DRAM[46311] = 8'b1111100;
DRAM[46312] = 8'b1111111;
DRAM[46313] = 8'b1111111;
DRAM[46314] = 8'b1111111;
DRAM[46315] = 8'b1111111;
DRAM[46316] = 8'b10000000;
DRAM[46317] = 8'b10000001;
DRAM[46318] = 8'b10000010;
DRAM[46319] = 8'b10000011;
DRAM[46320] = 8'b10000110;
DRAM[46321] = 8'b10000101;
DRAM[46322] = 8'b10000101;
DRAM[46323] = 8'b10000101;
DRAM[46324] = 8'b10000110;
DRAM[46325] = 8'b10001000;
DRAM[46326] = 8'b10001001;
DRAM[46327] = 8'b10001011;
DRAM[46328] = 8'b10001100;
DRAM[46329] = 8'b10001100;
DRAM[46330] = 8'b10001011;
DRAM[46331] = 8'b10001011;
DRAM[46332] = 8'b10001011;
DRAM[46333] = 8'b10001011;
DRAM[46334] = 8'b10001011;
DRAM[46335] = 8'b10001011;
DRAM[46336] = 8'b10001111;
DRAM[46337] = 8'b10001111;
DRAM[46338] = 8'b10001110;
DRAM[46339] = 8'b10001110;
DRAM[46340] = 8'b10001111;
DRAM[46341] = 8'b10010000;
DRAM[46342] = 8'b10010001;
DRAM[46343] = 8'b10010001;
DRAM[46344] = 8'b10010011;
DRAM[46345] = 8'b10010011;
DRAM[46346] = 8'b10010100;
DRAM[46347] = 8'b10010101;
DRAM[46348] = 8'b10010101;
DRAM[46349] = 8'b10010100;
DRAM[46350] = 8'b10010100;
DRAM[46351] = 8'b10010011;
DRAM[46352] = 8'b10010101;
DRAM[46353] = 8'b10010101;
DRAM[46354] = 8'b10010110;
DRAM[46355] = 8'b10010110;
DRAM[46356] = 8'b10010111;
DRAM[46357] = 8'b10011000;
DRAM[46358] = 8'b10011001;
DRAM[46359] = 8'b10011001;
DRAM[46360] = 8'b10011000;
DRAM[46361] = 8'b10011000;
DRAM[46362] = 8'b10011001;
DRAM[46363] = 8'b10011010;
DRAM[46364] = 8'b10011100;
DRAM[46365] = 8'b10100010;
DRAM[46366] = 8'b10101010;
DRAM[46367] = 8'b10101111;
DRAM[46368] = 8'b11001011;
DRAM[46369] = 8'b11011101;
DRAM[46370] = 8'b11110001;
DRAM[46371] = 8'b11111011;
DRAM[46372] = 8'b11111101;
DRAM[46373] = 8'b11111110;
DRAM[46374] = 8'b11111110;
DRAM[46375] = 8'b11111101;
DRAM[46376] = 8'b11111101;
DRAM[46377] = 8'b11111110;
DRAM[46378] = 8'b11111110;
DRAM[46379] = 8'b11111111;
DRAM[46380] = 8'b11111111;
DRAM[46381] = 8'b11111110;
DRAM[46382] = 8'b11111110;
DRAM[46383] = 8'b11111101;
DRAM[46384] = 8'b11111101;
DRAM[46385] = 8'b11111011;
DRAM[46386] = 8'b11111001;
DRAM[46387] = 8'b11111000;
DRAM[46388] = 8'b11111000;
DRAM[46389] = 8'b11110111;
DRAM[46390] = 8'b11110100;
DRAM[46391] = 8'b11110001;
DRAM[46392] = 8'b11110000;
DRAM[46393] = 8'b11101101;
DRAM[46394] = 8'b11101001;
DRAM[46395] = 8'b11100111;
DRAM[46396] = 8'b11100111;
DRAM[46397] = 8'b11101000;
DRAM[46398] = 8'b11100111;
DRAM[46399] = 8'b11100110;
DRAM[46400] = 8'b11100010;
DRAM[46401] = 8'b11011011;
DRAM[46402] = 8'b11010101;
DRAM[46403] = 8'b11010110;
DRAM[46404] = 8'b11011011;
DRAM[46405] = 8'b11011011;
DRAM[46406] = 8'b11010100;
DRAM[46407] = 8'b11001100;
DRAM[46408] = 8'b11000010;
DRAM[46409] = 8'b10111101;
DRAM[46410] = 8'b10110110;
DRAM[46411] = 8'b10110011;
DRAM[46412] = 8'b10110001;
DRAM[46413] = 8'b10101101;
DRAM[46414] = 8'b10101000;
DRAM[46415] = 8'b10100011;
DRAM[46416] = 8'b10100110;
DRAM[46417] = 8'b10101111;
DRAM[46418] = 8'b10110011;
DRAM[46419] = 8'b10101110;
DRAM[46420] = 8'b10101001;
DRAM[46421] = 8'b10100101;
DRAM[46422] = 8'b10011010;
DRAM[46423] = 8'b10001101;
DRAM[46424] = 8'b10010110;
DRAM[46425] = 8'b10001110;
DRAM[46426] = 8'b10000101;
DRAM[46427] = 8'b10000001;
DRAM[46428] = 8'b10000101;
DRAM[46429] = 8'b10001001;
DRAM[46430] = 8'b10001011;
DRAM[46431] = 8'b10001010;
DRAM[46432] = 8'b10000010;
DRAM[46433] = 8'b1111111;
DRAM[46434] = 8'b10000010;
DRAM[46435] = 8'b10001001;
DRAM[46436] = 8'b10001001;
DRAM[46437] = 8'b10000111;
DRAM[46438] = 8'b10001110;
DRAM[46439] = 8'b10011001;
DRAM[46440] = 8'b10100101;
DRAM[46441] = 8'b10011111;
DRAM[46442] = 8'b10011001;
DRAM[46443] = 8'b10010100;
DRAM[46444] = 8'b10001010;
DRAM[46445] = 8'b1111100;
DRAM[46446] = 8'b1110001;
DRAM[46447] = 8'b1101101;
DRAM[46448] = 8'b10011011;
DRAM[46449] = 8'b10101110;
DRAM[46450] = 8'b10111110;
DRAM[46451] = 8'b10111110;
DRAM[46452] = 8'b10110100;
DRAM[46453] = 8'b10101100;
DRAM[46454] = 8'b10101010;
DRAM[46455] = 8'b10101010;
DRAM[46456] = 8'b10011111;
DRAM[46457] = 8'b10100001;
DRAM[46458] = 8'b10011010;
DRAM[46459] = 8'b10001100;
DRAM[46460] = 8'b10000101;
DRAM[46461] = 8'b10000010;
DRAM[46462] = 8'b1111001;
DRAM[46463] = 8'b1101111;
DRAM[46464] = 8'b1101111;
DRAM[46465] = 8'b1100001;
DRAM[46466] = 8'b1001101;
DRAM[46467] = 8'b1000011;
DRAM[46468] = 8'b1000110;
DRAM[46469] = 8'b1001011;
DRAM[46470] = 8'b1000010;
DRAM[46471] = 8'b110100;
DRAM[46472] = 8'b110011;
DRAM[46473] = 8'b101001;
DRAM[46474] = 8'b11011;
DRAM[46475] = 8'b10011;
DRAM[46476] = 8'b10001;
DRAM[46477] = 8'b10011;
DRAM[46478] = 8'b10100;
DRAM[46479] = 8'b10100;
DRAM[46480] = 8'b11100;
DRAM[46481] = 8'b10101;
DRAM[46482] = 8'b10010;
DRAM[46483] = 8'b10011;
DRAM[46484] = 8'b1111;
DRAM[46485] = 8'b1000;
DRAM[46486] = 8'b1011;
DRAM[46487] = 8'b10011;
DRAM[46488] = 8'b11111;
DRAM[46489] = 8'b100011;
DRAM[46490] = 8'b100100;
DRAM[46491] = 8'b100001;
DRAM[46492] = 8'b100001;
DRAM[46493] = 8'b100100;
DRAM[46494] = 8'b100110;
DRAM[46495] = 8'b100101;
DRAM[46496] = 8'b101101;
DRAM[46497] = 8'b101100;
DRAM[46498] = 8'b101111;
DRAM[46499] = 8'b111000;
DRAM[46500] = 8'b1000100;
DRAM[46501] = 8'b1001111;
DRAM[46502] = 8'b1010110;
DRAM[46503] = 8'b1011010;
DRAM[46504] = 8'b1101100;
DRAM[46505] = 8'b1111010;
DRAM[46506] = 8'b10000110;
DRAM[46507] = 8'b10001100;
DRAM[46508] = 8'b10010110;
DRAM[46509] = 8'b10101000;
DRAM[46510] = 8'b10110110;
DRAM[46511] = 8'b10111011;
DRAM[46512] = 8'b11000110;
DRAM[46513] = 8'b11000110;
DRAM[46514] = 8'b11010001;
DRAM[46515] = 8'b11011100;
DRAM[46516] = 8'b11010100;
DRAM[46517] = 8'b11000100;
DRAM[46518] = 8'b11001011;
DRAM[46519] = 8'b11100000;
DRAM[46520] = 8'b11101100;
DRAM[46521] = 8'b11110011;
DRAM[46522] = 8'b11111010;
DRAM[46523] = 8'b11111101;
DRAM[46524] = 8'b11111101;
DRAM[46525] = 8'b11111101;
DRAM[46526] = 8'b11111110;
DRAM[46527] = 8'b11111111;
DRAM[46528] = 8'b11111110;
DRAM[46529] = 8'b11111011;
DRAM[46530] = 8'b11110101;
DRAM[46531] = 8'b11101011;
DRAM[46532] = 8'b11100011;
DRAM[46533] = 8'b11011010;
DRAM[46534] = 8'b11001101;
DRAM[46535] = 8'b11000001;
DRAM[46536] = 8'b10101110;
DRAM[46537] = 8'b10100110;
DRAM[46538] = 8'b10100001;
DRAM[46539] = 8'b10100010;
DRAM[46540] = 8'b10100010;
DRAM[46541] = 8'b10011101;
DRAM[46542] = 8'b10010111;
DRAM[46543] = 8'b10010011;
DRAM[46544] = 8'b10010110;
DRAM[46545] = 8'b10010011;
DRAM[46546] = 8'b10001110;
DRAM[46547] = 8'b10001010;
DRAM[46548] = 8'b10001001;
DRAM[46549] = 8'b10000111;
DRAM[46550] = 8'b10000110;
DRAM[46551] = 8'b10000100;
DRAM[46552] = 8'b10000101;
DRAM[46553] = 8'b10000011;
DRAM[46554] = 8'b10000000;
DRAM[46555] = 8'b10000000;
DRAM[46556] = 8'b10000000;
DRAM[46557] = 8'b10000001;
DRAM[46558] = 8'b10000000;
DRAM[46559] = 8'b1111110;
DRAM[46560] = 8'b1111100;
DRAM[46561] = 8'b1111100;
DRAM[46562] = 8'b1111100;
DRAM[46563] = 8'b1111100;
DRAM[46564] = 8'b1111100;
DRAM[46565] = 8'b1111100;
DRAM[46566] = 8'b1111100;
DRAM[46567] = 8'b1111100;
DRAM[46568] = 8'b10000000;
DRAM[46569] = 8'b10000000;
DRAM[46570] = 8'b10000000;
DRAM[46571] = 8'b10000000;
DRAM[46572] = 8'b10000000;
DRAM[46573] = 8'b10000001;
DRAM[46574] = 8'b10000010;
DRAM[46575] = 8'b10000011;
DRAM[46576] = 8'b10000110;
DRAM[46577] = 8'b10000101;
DRAM[46578] = 8'b10000101;
DRAM[46579] = 8'b10000101;
DRAM[46580] = 8'b10000110;
DRAM[46581] = 8'b10001000;
DRAM[46582] = 8'b10001010;
DRAM[46583] = 8'b10001100;
DRAM[46584] = 8'b10001101;
DRAM[46585] = 8'b10001101;
DRAM[46586] = 8'b10001100;
DRAM[46587] = 8'b10001011;
DRAM[46588] = 8'b10001011;
DRAM[46589] = 8'b10001011;
DRAM[46590] = 8'b10001011;
DRAM[46591] = 8'b10001100;
DRAM[46592] = 8'b10001111;
DRAM[46593] = 8'b10001111;
DRAM[46594] = 8'b10001110;
DRAM[46595] = 8'b10001110;
DRAM[46596] = 8'b10001111;
DRAM[46597] = 8'b10001111;
DRAM[46598] = 8'b10010000;
DRAM[46599] = 8'b10010001;
DRAM[46600] = 8'b10001111;
DRAM[46601] = 8'b10001111;
DRAM[46602] = 8'b10010001;
DRAM[46603] = 8'b10010010;
DRAM[46604] = 8'b10010010;
DRAM[46605] = 8'b10010010;
DRAM[46606] = 8'b10010010;
DRAM[46607] = 8'b10010010;
DRAM[46608] = 8'b10010100;
DRAM[46609] = 8'b10010100;
DRAM[46610] = 8'b10010101;
DRAM[46611] = 8'b10010110;
DRAM[46612] = 8'b10010111;
DRAM[46613] = 8'b10010111;
DRAM[46614] = 8'b10011000;
DRAM[46615] = 8'b10011000;
DRAM[46616] = 8'b10010111;
DRAM[46617] = 8'b10011000;
DRAM[46618] = 8'b10011010;
DRAM[46619] = 8'b10011011;
DRAM[46620] = 8'b10011110;
DRAM[46621] = 8'b10100110;
DRAM[46622] = 8'b10101111;
DRAM[46623] = 8'b10110111;
DRAM[46624] = 8'b11010100;
DRAM[46625] = 8'b11100100;
DRAM[46626] = 8'b11110100;
DRAM[46627] = 8'b11111001;
DRAM[46628] = 8'b11111011;
DRAM[46629] = 8'b11111110;
DRAM[46630] = 8'b11111111;
DRAM[46631] = 8'b11111110;
DRAM[46632] = 8'b11111101;
DRAM[46633] = 8'b11111110;
DRAM[46634] = 8'b11111110;
DRAM[46635] = 8'b11111111;
DRAM[46636] = 8'b11111111;
DRAM[46637] = 8'b11111110;
DRAM[46638] = 8'b11111110;
DRAM[46639] = 8'b11111101;
DRAM[46640] = 8'b11111110;
DRAM[46641] = 8'b11111100;
DRAM[46642] = 8'b11111001;
DRAM[46643] = 8'b11110111;
DRAM[46644] = 8'b11110111;
DRAM[46645] = 8'b11110111;
DRAM[46646] = 8'b11110110;
DRAM[46647] = 8'b11110101;
DRAM[46648] = 8'b11101110;
DRAM[46649] = 8'b11101101;
DRAM[46650] = 8'b11101011;
DRAM[46651] = 8'b11101011;
DRAM[46652] = 8'b11101100;
DRAM[46653] = 8'b11101100;
DRAM[46654] = 8'b11101010;
DRAM[46655] = 8'b11101000;
DRAM[46656] = 8'b11101000;
DRAM[46657] = 8'b11011111;
DRAM[46658] = 8'b11010110;
DRAM[46659] = 8'b11010100;
DRAM[46660] = 8'b11010101;
DRAM[46661] = 8'b11010010;
DRAM[46662] = 8'b11001001;
DRAM[46663] = 8'b11000000;
DRAM[46664] = 8'b11001000;
DRAM[46665] = 8'b11000010;
DRAM[46666] = 8'b10111011;
DRAM[46667] = 8'b10110101;
DRAM[46668] = 8'b10110011;
DRAM[46669] = 8'b10101111;
DRAM[46670] = 8'b10100111;
DRAM[46671] = 8'b10011111;
DRAM[46672] = 8'b10100010;
DRAM[46673] = 8'b10110010;
DRAM[46674] = 8'b10110111;
DRAM[46675] = 8'b10101000;
DRAM[46676] = 8'b10011001;
DRAM[46677] = 8'b10010111;
DRAM[46678] = 8'b10011100;
DRAM[46679] = 8'b10011101;
DRAM[46680] = 8'b10010011;
DRAM[46681] = 8'b10001101;
DRAM[46682] = 8'b10000111;
DRAM[46683] = 8'b10000111;
DRAM[46684] = 8'b10001010;
DRAM[46685] = 8'b10001100;
DRAM[46686] = 8'b10001001;
DRAM[46687] = 8'b10000110;
DRAM[46688] = 8'b10001101;
DRAM[46689] = 8'b10001001;
DRAM[46690] = 8'b10001001;
DRAM[46691] = 8'b10001100;
DRAM[46692] = 8'b10000111;
DRAM[46693] = 8'b1111111;
DRAM[46694] = 8'b10000010;
DRAM[46695] = 8'b10001101;
DRAM[46696] = 8'b10011100;
DRAM[46697] = 8'b10101001;
DRAM[46698] = 8'b10101100;
DRAM[46699] = 8'b10010111;
DRAM[46700] = 8'b1111100;
DRAM[46701] = 8'b1110000;
DRAM[46702] = 8'b1111000;
DRAM[46703] = 8'b10000100;
DRAM[46704] = 8'b10001000;
DRAM[46705] = 8'b10011110;
DRAM[46706] = 8'b10110011;
DRAM[46707] = 8'b10110110;
DRAM[46708] = 8'b10101101;
DRAM[46709] = 8'b10100111;
DRAM[46710] = 8'b10101001;
DRAM[46711] = 8'b10101100;
DRAM[46712] = 8'b10101000;
DRAM[46713] = 8'b10101010;
DRAM[46714] = 8'b10100000;
DRAM[46715] = 8'b10010010;
DRAM[46716] = 8'b10000110;
DRAM[46717] = 8'b1110110;
DRAM[46718] = 8'b1101001;
DRAM[46719] = 8'b1101000;
DRAM[46720] = 8'b1101101;
DRAM[46721] = 8'b1011110;
DRAM[46722] = 8'b1001100;
DRAM[46723] = 8'b1001000;
DRAM[46724] = 8'b1010000;
DRAM[46725] = 8'b1010010;
DRAM[46726] = 8'b1000100;
DRAM[46727] = 8'b110001;
DRAM[46728] = 8'b110110;
DRAM[46729] = 8'b101010;
DRAM[46730] = 8'b11101;
DRAM[46731] = 8'b11000;
DRAM[46732] = 8'b11100;
DRAM[46733] = 8'b100001;
DRAM[46734] = 8'b100001;
DRAM[46735] = 8'b11110;
DRAM[46736] = 8'b101000;
DRAM[46737] = 8'b11101;
DRAM[46738] = 8'b10110;
DRAM[46739] = 8'b10100;
DRAM[46740] = 8'b1101;
DRAM[46741] = 8'b101;
DRAM[46742] = 8'b1000;
DRAM[46743] = 8'b10010;
DRAM[46744] = 8'b11001;
DRAM[46745] = 8'b11110;
DRAM[46746] = 8'b100011;
DRAM[46747] = 8'b100110;
DRAM[46748] = 8'b101100;
DRAM[46749] = 8'b110001;
DRAM[46750] = 8'b101111;
DRAM[46751] = 8'b101011;
DRAM[46752] = 8'b101111;
DRAM[46753] = 8'b110000;
DRAM[46754] = 8'b110010;
DRAM[46755] = 8'b110101;
DRAM[46756] = 8'b111101;
DRAM[46757] = 8'b1001000;
DRAM[46758] = 8'b1010001;
DRAM[46759] = 8'b1010110;
DRAM[46760] = 8'b1011100;
DRAM[46761] = 8'b1101111;
DRAM[46762] = 8'b1111110;
DRAM[46763] = 8'b10000101;
DRAM[46764] = 8'b10010000;
DRAM[46765] = 8'b10100010;
DRAM[46766] = 8'b10101101;
DRAM[46767] = 8'b10101100;
DRAM[46768] = 8'b11000010;
DRAM[46769] = 8'b11010100;
DRAM[46770] = 8'b11011011;
DRAM[46771] = 8'b11010000;
DRAM[46772] = 8'b11001001;
DRAM[46773] = 8'b11010010;
DRAM[46774] = 8'b11100010;
DRAM[46775] = 8'b11101010;
DRAM[46776] = 8'b11110011;
DRAM[46777] = 8'b11110110;
DRAM[46778] = 8'b11111010;
DRAM[46779] = 8'b11111101;
DRAM[46780] = 8'b11111100;
DRAM[46781] = 8'b11111100;
DRAM[46782] = 8'b11111110;
DRAM[46783] = 8'b11111111;
DRAM[46784] = 8'b11111010;
DRAM[46785] = 8'b11111010;
DRAM[46786] = 8'b11110011;
DRAM[46787] = 8'b11100110;
DRAM[46788] = 8'b11011010;
DRAM[46789] = 8'b11010010;
DRAM[46790] = 8'b11001000;
DRAM[46791] = 8'b10111110;
DRAM[46792] = 8'b10101111;
DRAM[46793] = 8'b10101100;
DRAM[46794] = 8'b10100101;
DRAM[46795] = 8'b10011110;
DRAM[46796] = 8'b10011100;
DRAM[46797] = 8'b10011100;
DRAM[46798] = 8'b10011000;
DRAM[46799] = 8'b10010001;
DRAM[46800] = 8'b10011000;
DRAM[46801] = 8'b10010011;
DRAM[46802] = 8'b10001100;
DRAM[46803] = 8'b10000111;
DRAM[46804] = 8'b10000110;
DRAM[46805] = 8'b10000101;
DRAM[46806] = 8'b10000101;
DRAM[46807] = 8'b10000100;
DRAM[46808] = 8'b10000011;
DRAM[46809] = 8'b10000001;
DRAM[46810] = 8'b1111110;
DRAM[46811] = 8'b1111110;
DRAM[46812] = 8'b1111110;
DRAM[46813] = 8'b1111111;
DRAM[46814] = 8'b1111110;
DRAM[46815] = 8'b1111100;
DRAM[46816] = 8'b1111011;
DRAM[46817] = 8'b1111011;
DRAM[46818] = 8'b1111011;
DRAM[46819] = 8'b1111011;
DRAM[46820] = 8'b1111011;
DRAM[46821] = 8'b1111011;
DRAM[46822] = 8'b1111011;
DRAM[46823] = 8'b1111011;
DRAM[46824] = 8'b10000001;
DRAM[46825] = 8'b10000000;
DRAM[46826] = 8'b10000000;
DRAM[46827] = 8'b10000000;
DRAM[46828] = 8'b10000000;
DRAM[46829] = 8'b10000001;
DRAM[46830] = 8'b10000010;
DRAM[46831] = 8'b10000011;
DRAM[46832] = 8'b10000110;
DRAM[46833] = 8'b10000101;
DRAM[46834] = 8'b10000100;
DRAM[46835] = 8'b10000100;
DRAM[46836] = 8'b10000101;
DRAM[46837] = 8'b10001000;
DRAM[46838] = 8'b10001011;
DRAM[46839] = 8'b10001100;
DRAM[46840] = 8'b10001110;
DRAM[46841] = 8'b10001101;
DRAM[46842] = 8'b10001100;
DRAM[46843] = 8'b10001011;
DRAM[46844] = 8'b10001010;
DRAM[46845] = 8'b10001011;
DRAM[46846] = 8'b10001011;
DRAM[46847] = 8'b10001100;
DRAM[46848] = 8'b10001111;
DRAM[46849] = 8'b10001110;
DRAM[46850] = 8'b10001110;
DRAM[46851] = 8'b10001110;
DRAM[46852] = 8'b10001110;
DRAM[46853] = 8'b10001111;
DRAM[46854] = 8'b10010000;
DRAM[46855] = 8'b10010001;
DRAM[46856] = 8'b10001011;
DRAM[46857] = 8'b10001100;
DRAM[46858] = 8'b10001110;
DRAM[46859] = 8'b10001111;
DRAM[46860] = 8'b10010000;
DRAM[46861] = 8'b10010001;
DRAM[46862] = 8'b10010001;
DRAM[46863] = 8'b10010001;
DRAM[46864] = 8'b10010100;
DRAM[46865] = 8'b10010100;
DRAM[46866] = 8'b10010101;
DRAM[46867] = 8'b10010101;
DRAM[46868] = 8'b10010110;
DRAM[46869] = 8'b10010111;
DRAM[46870] = 8'b10011000;
DRAM[46871] = 8'b10011000;
DRAM[46872] = 8'b10010111;
DRAM[46873] = 8'b10011001;
DRAM[46874] = 8'b10011010;
DRAM[46875] = 8'b10011100;
DRAM[46876] = 8'b10100000;
DRAM[46877] = 8'b10101000;
DRAM[46878] = 8'b10110011;
DRAM[46879] = 8'b10111011;
DRAM[46880] = 8'b11010110;
DRAM[46881] = 8'b11100101;
DRAM[46882] = 8'b11110001;
DRAM[46883] = 8'b11110101;
DRAM[46884] = 8'b11111000;
DRAM[46885] = 8'b11111101;
DRAM[46886] = 8'b11111111;
DRAM[46887] = 8'b11111101;
DRAM[46888] = 8'b11111101;
DRAM[46889] = 8'b11111110;
DRAM[46890] = 8'b11111110;
DRAM[46891] = 8'b11111111;
DRAM[46892] = 8'b11111111;
DRAM[46893] = 8'b11111110;
DRAM[46894] = 8'b11111110;
DRAM[46895] = 8'b11111101;
DRAM[46896] = 8'b11111010;
DRAM[46897] = 8'b11110111;
DRAM[46898] = 8'b11110011;
DRAM[46899] = 8'b11110001;
DRAM[46900] = 8'b11110010;
DRAM[46901] = 8'b11110011;
DRAM[46902] = 8'b11110011;
DRAM[46903] = 8'b11110010;
DRAM[46904] = 8'b11110000;
DRAM[46905] = 8'b11101111;
DRAM[46906] = 8'b11101111;
DRAM[46907] = 8'b11101111;
DRAM[46908] = 8'b11101110;
DRAM[46909] = 8'b11101011;
DRAM[46910] = 8'b11100110;
DRAM[46911] = 8'b11100001;
DRAM[46912] = 8'b11010111;
DRAM[46913] = 8'b11011010;
DRAM[46914] = 8'b11011011;
DRAM[46915] = 8'b11010111;
DRAM[46916] = 8'b11001111;
DRAM[46917] = 8'b11001010;
DRAM[46918] = 8'b11001001;
DRAM[46919] = 8'b11001011;
DRAM[46920] = 8'b11000010;
DRAM[46921] = 8'b11000000;
DRAM[46922] = 8'b10111101;
DRAM[46923] = 8'b10111100;
DRAM[46924] = 8'b10111011;
DRAM[46925] = 8'b10110110;
DRAM[46926] = 8'b10101001;
DRAM[46927] = 8'b10011101;
DRAM[46928] = 8'b10101101;
DRAM[46929] = 8'b10101101;
DRAM[46930] = 8'b10100100;
DRAM[46931] = 8'b10010111;
DRAM[46932] = 8'b10010111;
DRAM[46933] = 8'b10100010;
DRAM[46934] = 8'b10100110;
DRAM[46935] = 8'b10100000;
DRAM[46936] = 8'b10010111;
DRAM[46937] = 8'b10010101;
DRAM[46938] = 8'b10010100;
DRAM[46939] = 8'b10010101;
DRAM[46940] = 8'b10010101;
DRAM[46941] = 8'b10010011;
DRAM[46942] = 8'b10001110;
DRAM[46943] = 8'b10001010;
DRAM[46944] = 8'b10001001;
DRAM[46945] = 8'b10000100;
DRAM[46946] = 8'b10000100;
DRAM[46947] = 8'b10001000;
DRAM[46948] = 8'b10000101;
DRAM[46949] = 8'b1111111;
DRAM[46950] = 8'b10000110;
DRAM[46951] = 8'b10010100;
DRAM[46952] = 8'b10010111;
DRAM[46953] = 8'b10100001;
DRAM[46954] = 8'b10100011;
DRAM[46955] = 8'b10010111;
DRAM[46956] = 8'b10001110;
DRAM[46957] = 8'b10001110;
DRAM[46958] = 8'b10001100;
DRAM[46959] = 8'b10000110;
DRAM[46960] = 8'b10000001;
DRAM[46961] = 8'b10010000;
DRAM[46962] = 8'b10100000;
DRAM[46963] = 8'b10101001;
DRAM[46964] = 8'b10101110;
DRAM[46965] = 8'b10110000;
DRAM[46966] = 8'b10101110;
DRAM[46967] = 8'b10101010;
DRAM[46968] = 8'b10100101;
DRAM[46969] = 8'b10100111;
DRAM[46970] = 8'b10100000;
DRAM[46971] = 8'b10010101;
DRAM[46972] = 8'b10001011;
DRAM[46973] = 8'b1110111;
DRAM[46974] = 8'b1101011;
DRAM[46975] = 8'b1110010;
DRAM[46976] = 8'b1101000;
DRAM[46977] = 8'b1100011;
DRAM[46978] = 8'b1011101;
DRAM[46979] = 8'b1011001;
DRAM[46980] = 8'b1011001;
DRAM[46981] = 8'b1010011;
DRAM[46982] = 8'b1000110;
DRAM[46983] = 8'b111001;
DRAM[46984] = 8'b110010;
DRAM[46985] = 8'b100110;
DRAM[46986] = 8'b11011;
DRAM[46987] = 8'b11010;
DRAM[46988] = 8'b100011;
DRAM[46989] = 8'b101010;
DRAM[46990] = 8'b101000;
DRAM[46991] = 8'b100011;
DRAM[46992] = 8'b101000;
DRAM[46993] = 8'b11010;
DRAM[46994] = 8'b1111;
DRAM[46995] = 8'b1010;
DRAM[46996] = 8'b10;
DRAM[46997] = 8'b0;
DRAM[46998] = 8'b0;
DRAM[46999] = 8'b1010;
DRAM[47000] = 8'b111;
DRAM[47001] = 8'b1110;
DRAM[47002] = 8'b10111;
DRAM[47003] = 8'b100000;
DRAM[47004] = 8'b101010;
DRAM[47005] = 8'b110000;
DRAM[47006] = 8'b101100;
DRAM[47007] = 8'b100100;
DRAM[47008] = 8'b110010;
DRAM[47009] = 8'b110110;
DRAM[47010] = 8'b111000;
DRAM[47011] = 8'b110111;
DRAM[47012] = 8'b111001;
DRAM[47013] = 8'b1000011;
DRAM[47014] = 8'b1010000;
DRAM[47015] = 8'b1011000;
DRAM[47016] = 8'b1010101;
DRAM[47017] = 8'b1101001;
DRAM[47018] = 8'b1111010;
DRAM[47019] = 8'b10000010;
DRAM[47020] = 8'b10010001;
DRAM[47021] = 8'b10100101;
DRAM[47022] = 8'b10101100;
DRAM[47023] = 8'b10100111;
DRAM[47024] = 8'b11000110;
DRAM[47025] = 8'b11100101;
DRAM[47026] = 8'b11100111;
DRAM[47027] = 8'b11000101;
DRAM[47028] = 8'b10111100;
DRAM[47029] = 8'b11011010;
DRAM[47030] = 8'b11101110;
DRAM[47031] = 8'b11101000;
DRAM[47032] = 8'b11110110;
DRAM[47033] = 8'b11110111;
DRAM[47034] = 8'b11111010;
DRAM[47035] = 8'b11111100;
DRAM[47036] = 8'b11111100;
DRAM[47037] = 8'b11111011;
DRAM[47038] = 8'b11111110;
DRAM[47039] = 8'b11111111;
DRAM[47040] = 8'b11111100;
DRAM[47041] = 8'b11111101;
DRAM[47042] = 8'b11110110;
DRAM[47043] = 8'b11100110;
DRAM[47044] = 8'b11010111;
DRAM[47045] = 8'b11001111;
DRAM[47046] = 8'b11000111;
DRAM[47047] = 8'b10111110;
DRAM[47048] = 8'b10101111;
DRAM[47049] = 8'b10110001;
DRAM[47050] = 8'b10101001;
DRAM[47051] = 8'b10011011;
DRAM[47052] = 8'b10010101;
DRAM[47053] = 8'b10011001;
DRAM[47054] = 8'b10011001;
DRAM[47055] = 8'b10010011;
DRAM[47056] = 8'b10011000;
DRAM[47057] = 8'b10010010;
DRAM[47058] = 8'b10001010;
DRAM[47059] = 8'b10000101;
DRAM[47060] = 8'b10000011;
DRAM[47061] = 8'b10000011;
DRAM[47062] = 8'b10000100;
DRAM[47063] = 8'b10000100;
DRAM[47064] = 8'b10000001;
DRAM[47065] = 8'b1111111;
DRAM[47066] = 8'b1111100;
DRAM[47067] = 8'b1111100;
DRAM[47068] = 8'b1111100;
DRAM[47069] = 8'b1111101;
DRAM[47070] = 8'b1111100;
DRAM[47071] = 8'b1111010;
DRAM[47072] = 8'b1111011;
DRAM[47073] = 8'b1111011;
DRAM[47074] = 8'b1111011;
DRAM[47075] = 8'b1111011;
DRAM[47076] = 8'b1111011;
DRAM[47077] = 8'b1111011;
DRAM[47078] = 8'b1111011;
DRAM[47079] = 8'b1111011;
DRAM[47080] = 8'b10000001;
DRAM[47081] = 8'b10000001;
DRAM[47082] = 8'b10000000;
DRAM[47083] = 8'b10000000;
DRAM[47084] = 8'b10000000;
DRAM[47085] = 8'b10000001;
DRAM[47086] = 8'b10000010;
DRAM[47087] = 8'b10000010;
DRAM[47088] = 8'b10000110;
DRAM[47089] = 8'b10000101;
DRAM[47090] = 8'b10000100;
DRAM[47091] = 8'b10000100;
DRAM[47092] = 8'b10000101;
DRAM[47093] = 8'b10001000;
DRAM[47094] = 8'b10001011;
DRAM[47095] = 8'b10001101;
DRAM[47096] = 8'b10001111;
DRAM[47097] = 8'b10001110;
DRAM[47098] = 8'b10001100;
DRAM[47099] = 8'b10001011;
DRAM[47100] = 8'b10001010;
DRAM[47101] = 8'b10001011;
DRAM[47102] = 8'b10001011;
DRAM[47103] = 8'b10001100;
DRAM[47104] = 8'b10001110;
DRAM[47105] = 8'b10001100;
DRAM[47106] = 8'b10001100;
DRAM[47107] = 8'b10001100;
DRAM[47108] = 8'b10001110;
DRAM[47109] = 8'b10001111;
DRAM[47110] = 8'b10001110;
DRAM[47111] = 8'b10001101;
DRAM[47112] = 8'b10001110;
DRAM[47113] = 8'b10001111;
DRAM[47114] = 8'b10001111;
DRAM[47115] = 8'b10010001;
DRAM[47116] = 8'b10010010;
DRAM[47117] = 8'b10010011;
DRAM[47118] = 8'b10010100;
DRAM[47119] = 8'b10010100;
DRAM[47120] = 8'b10010100;
DRAM[47121] = 8'b10010100;
DRAM[47122] = 8'b10010101;
DRAM[47123] = 8'b10010101;
DRAM[47124] = 8'b10010101;
DRAM[47125] = 8'b10010110;
DRAM[47126] = 8'b10010110;
DRAM[47127] = 8'b10010110;
DRAM[47128] = 8'b10011010;
DRAM[47129] = 8'b10011100;
DRAM[47130] = 8'b10011000;
DRAM[47131] = 8'b10011011;
DRAM[47132] = 8'b10100111;
DRAM[47133] = 8'b10101011;
DRAM[47134] = 8'b10110001;
DRAM[47135] = 8'b11000000;
DRAM[47136] = 8'b11001011;
DRAM[47137] = 8'b11001111;
DRAM[47138] = 8'b11011100;
DRAM[47139] = 8'b11101111;
DRAM[47140] = 8'b11111110;
DRAM[47141] = 8'b11111111;
DRAM[47142] = 8'b11111111;
DRAM[47143] = 8'b11111011;
DRAM[47144] = 8'b11111111;
DRAM[47145] = 8'b11111111;
DRAM[47146] = 8'b11111110;
DRAM[47147] = 8'b11111101;
DRAM[47148] = 8'b11111101;
DRAM[47149] = 8'b11111101;
DRAM[47150] = 8'b11111110;
DRAM[47151] = 8'b11111110;
DRAM[47152] = 8'b11110111;
DRAM[47153] = 8'b11111001;
DRAM[47154] = 8'b11111011;
DRAM[47155] = 8'b11111011;
DRAM[47156] = 8'b11111000;
DRAM[47157] = 8'b11110100;
DRAM[47158] = 8'b11110001;
DRAM[47159] = 8'b11101111;
DRAM[47160] = 8'b11110010;
DRAM[47161] = 8'b11110001;
DRAM[47162] = 8'b11101101;
DRAM[47163] = 8'b11101001;
DRAM[47164] = 8'b11100100;
DRAM[47165] = 8'b11100001;
DRAM[47166] = 8'b11100000;
DRAM[47167] = 8'b11100001;
DRAM[47168] = 8'b11011000;
DRAM[47169] = 8'b11010100;
DRAM[47170] = 8'b11010010;
DRAM[47171] = 8'b11010011;
DRAM[47172] = 8'b11001110;
DRAM[47173] = 8'b11000101;
DRAM[47174] = 8'b11000011;
DRAM[47175] = 8'b11000111;
DRAM[47176] = 8'b11000001;
DRAM[47177] = 8'b10111110;
DRAM[47178] = 8'b10111111;
DRAM[47179] = 8'b11000000;
DRAM[47180] = 8'b10111011;
DRAM[47181] = 8'b10110011;
DRAM[47182] = 8'b10110010;
DRAM[47183] = 8'b10110110;
DRAM[47184] = 8'b10101000;
DRAM[47185] = 8'b10100010;
DRAM[47186] = 8'b10010110;
DRAM[47187] = 8'b10001111;
DRAM[47188] = 8'b10011000;
DRAM[47189] = 8'b10100110;
DRAM[47190] = 8'b10100101;
DRAM[47191] = 8'b10011010;
DRAM[47192] = 8'b10100000;
DRAM[47193] = 8'b10011111;
DRAM[47194] = 8'b10010101;
DRAM[47195] = 8'b10010001;
DRAM[47196] = 8'b10010111;
DRAM[47197] = 8'b10010001;
DRAM[47198] = 8'b10000111;
DRAM[47199] = 8'b10001001;
DRAM[47200] = 8'b1110000;
DRAM[47201] = 8'b1111101;
DRAM[47202] = 8'b1111111;
DRAM[47203] = 8'b1111001;
DRAM[47204] = 8'b1111110;
DRAM[47205] = 8'b10010000;
DRAM[47206] = 8'b10010111;
DRAM[47207] = 8'b10010001;
DRAM[47208] = 8'b10001100;
DRAM[47209] = 8'b10010110;
DRAM[47210] = 8'b10011111;
DRAM[47211] = 8'b10011110;
DRAM[47212] = 8'b10011001;
DRAM[47213] = 8'b10010100;
DRAM[47214] = 8'b10001110;
DRAM[47215] = 8'b10001001;
DRAM[47216] = 8'b1110010;
DRAM[47217] = 8'b1101100;
DRAM[47218] = 8'b1111010;
DRAM[47219] = 8'b10011100;
DRAM[47220] = 8'b10110010;
DRAM[47221] = 8'b10101101;
DRAM[47222] = 8'b10100011;
DRAM[47223] = 8'b10100000;
DRAM[47224] = 8'b10011101;
DRAM[47225] = 8'b10100110;
DRAM[47226] = 8'b10011011;
DRAM[47227] = 8'b1111111;
DRAM[47228] = 8'b1110011;
DRAM[47229] = 8'b1111010;
DRAM[47230] = 8'b1110101;
DRAM[47231] = 8'b1100100;
DRAM[47232] = 8'b1100110;
DRAM[47233] = 8'b1100000;
DRAM[47234] = 8'b1011000;
DRAM[47235] = 8'b1010011;
DRAM[47236] = 8'b1010010;
DRAM[47237] = 8'b1001101;
DRAM[47238] = 8'b1000000;
DRAM[47239] = 8'b110011;
DRAM[47240] = 8'b101010;
DRAM[47241] = 8'b100101;
DRAM[47242] = 8'b100011;
DRAM[47243] = 8'b101001;
DRAM[47244] = 8'b101110;
DRAM[47245] = 8'b101100;
DRAM[47246] = 8'b100101;
DRAM[47247] = 8'b11111;
DRAM[47248] = 8'b10011;
DRAM[47249] = 8'b1111;
DRAM[47250] = 8'b111;
DRAM[47251] = 8'b0;
DRAM[47252] = 8'b0;
DRAM[47253] = 8'b0;
DRAM[47254] = 8'b10;
DRAM[47255] = 8'b10;
DRAM[47256] = 8'b1000;
DRAM[47257] = 8'b111;
DRAM[47258] = 8'b101;
DRAM[47259] = 8'b1101;
DRAM[47260] = 8'b10110;
DRAM[47261] = 8'b1111;
DRAM[47262] = 8'b1110;
DRAM[47263] = 8'b11100;
DRAM[47264] = 8'b11111;
DRAM[47265] = 8'b101011;
DRAM[47266] = 8'b101111;
DRAM[47267] = 8'b110101;
DRAM[47268] = 8'b1000110;
DRAM[47269] = 8'b1010000;
DRAM[47270] = 8'b1010101;
DRAM[47271] = 8'b1011110;
DRAM[47272] = 8'b1011110;
DRAM[47273] = 8'b1101011;
DRAM[47274] = 8'b1111110;
DRAM[47275] = 8'b10001101;
DRAM[47276] = 8'b10010110;
DRAM[47277] = 8'b10011111;
DRAM[47278] = 8'b10101111;
DRAM[47279] = 8'b10111101;
DRAM[47280] = 8'b11010010;
DRAM[47281] = 8'b11001111;
DRAM[47282] = 8'b11001010;
DRAM[47283] = 8'b11000111;
DRAM[47284] = 8'b11001001;
DRAM[47285] = 8'b11010011;
DRAM[47286] = 8'b11100001;
DRAM[47287] = 8'b11101100;
DRAM[47288] = 8'b11110010;
DRAM[47289] = 8'b11110101;
DRAM[47290] = 8'b11111001;
DRAM[47291] = 8'b11111100;
DRAM[47292] = 8'b11111110;
DRAM[47293] = 8'b11111110;
DRAM[47294] = 8'b11111101;
DRAM[47295] = 8'b11111011;
DRAM[47296] = 8'b11111110;
DRAM[47297] = 8'b11111010;
DRAM[47298] = 8'b11110001;
DRAM[47299] = 8'b11100100;
DRAM[47300] = 8'b11010101;
DRAM[47301] = 8'b11001011;
DRAM[47302] = 8'b11000110;
DRAM[47303] = 8'b11000100;
DRAM[47304] = 8'b10110100;
DRAM[47305] = 8'b10101000;
DRAM[47306] = 8'b10100100;
DRAM[47307] = 8'b10101001;
DRAM[47308] = 8'b10100100;
DRAM[47309] = 8'b10010100;
DRAM[47310] = 8'b10001110;
DRAM[47311] = 8'b10010011;
DRAM[47312] = 8'b10001100;
DRAM[47313] = 8'b10001010;
DRAM[47314] = 8'b10000110;
DRAM[47315] = 8'b10000100;
DRAM[47316] = 8'b10000011;
DRAM[47317] = 8'b10000010;
DRAM[47318] = 8'b10000000;
DRAM[47319] = 8'b1111110;
DRAM[47320] = 8'b1111100;
DRAM[47321] = 8'b1111101;
DRAM[47322] = 8'b1111110;
DRAM[47323] = 8'b1111110;
DRAM[47324] = 8'b1111110;
DRAM[47325] = 8'b1111100;
DRAM[47326] = 8'b1111010;
DRAM[47327] = 8'b1111001;
DRAM[47328] = 8'b1111000;
DRAM[47329] = 8'b1111000;
DRAM[47330] = 8'b1111001;
DRAM[47331] = 8'b1111010;
DRAM[47332] = 8'b1111010;
DRAM[47333] = 8'b1111011;
DRAM[47334] = 8'b1111100;
DRAM[47335] = 8'b1111100;
DRAM[47336] = 8'b10000010;
DRAM[47337] = 8'b10000001;
DRAM[47338] = 8'b10000000;
DRAM[47339] = 8'b1111101;
DRAM[47340] = 8'b1111100;
DRAM[47341] = 8'b1111110;
DRAM[47342] = 8'b10000010;
DRAM[47343] = 8'b10000101;
DRAM[47344] = 8'b10000010;
DRAM[47345] = 8'b10000011;
DRAM[47346] = 8'b10000011;
DRAM[47347] = 8'b10000100;
DRAM[47348] = 8'b10000110;
DRAM[47349] = 8'b10001000;
DRAM[47350] = 8'b10001010;
DRAM[47351] = 8'b10001011;
DRAM[47352] = 8'b10001011;
DRAM[47353] = 8'b10001011;
DRAM[47354] = 8'b10001011;
DRAM[47355] = 8'b10001010;
DRAM[47356] = 8'b10001010;
DRAM[47357] = 8'b10001001;
DRAM[47358] = 8'b10001001;
DRAM[47359] = 8'b10001001;
DRAM[47360] = 8'b10001011;
DRAM[47361] = 8'b10001001;
DRAM[47362] = 8'b10001000;
DRAM[47363] = 8'b10001001;
DRAM[47364] = 8'b10001011;
DRAM[47365] = 8'b10001100;
DRAM[47366] = 8'b10001011;
DRAM[47367] = 8'b10001010;
DRAM[47368] = 8'b10001101;
DRAM[47369] = 8'b10001101;
DRAM[47370] = 8'b10001110;
DRAM[47371] = 8'b10001111;
DRAM[47372] = 8'b10010001;
DRAM[47373] = 8'b10010010;
DRAM[47374] = 8'b10010011;
DRAM[47375] = 8'b10010011;
DRAM[47376] = 8'b10010011;
DRAM[47377] = 8'b10010011;
DRAM[47378] = 8'b10010100;
DRAM[47379] = 8'b10010100;
DRAM[47380] = 8'b10010101;
DRAM[47381] = 8'b10010101;
DRAM[47382] = 8'b10010110;
DRAM[47383] = 8'b10010110;
DRAM[47384] = 8'b10011001;
DRAM[47385] = 8'b10011100;
DRAM[47386] = 8'b10011000;
DRAM[47387] = 8'b10011011;
DRAM[47388] = 8'b10100110;
DRAM[47389] = 8'b10101000;
DRAM[47390] = 8'b10101100;
DRAM[47391] = 8'b10111010;
DRAM[47392] = 8'b10111011;
DRAM[47393] = 8'b11001000;
DRAM[47394] = 8'b11011101;
DRAM[47395] = 8'b11110000;
DRAM[47396] = 8'b11111011;
DRAM[47397] = 8'b11111101;
DRAM[47398] = 8'b11111100;
DRAM[47399] = 8'b11111100;
DRAM[47400] = 8'b11111110;
DRAM[47401] = 8'b11111110;
DRAM[47402] = 8'b11111101;
DRAM[47403] = 8'b11111101;
DRAM[47404] = 8'b11111100;
DRAM[47405] = 8'b11111101;
DRAM[47406] = 8'b11111101;
DRAM[47407] = 8'b11111101;
DRAM[47408] = 8'b11111101;
DRAM[47409] = 8'b11111100;
DRAM[47410] = 8'b11111001;
DRAM[47411] = 8'b11110110;
DRAM[47412] = 8'b11110010;
DRAM[47413] = 8'b11101111;
DRAM[47414] = 8'b11101110;
DRAM[47415] = 8'b11101101;
DRAM[47416] = 8'b11100111;
DRAM[47417] = 8'b11100101;
DRAM[47418] = 8'b11100010;
DRAM[47419] = 8'b11011110;
DRAM[47420] = 8'b11011011;
DRAM[47421] = 8'b11011001;
DRAM[47422] = 8'b11011000;
DRAM[47423] = 8'b11011001;
DRAM[47424] = 8'b11010010;
DRAM[47425] = 8'b11001111;
DRAM[47426] = 8'b11001111;
DRAM[47427] = 8'b11001111;
DRAM[47428] = 8'b11001001;
DRAM[47429] = 8'b11000010;
DRAM[47430] = 8'b11000011;
DRAM[47431] = 8'b11001000;
DRAM[47432] = 8'b10111101;
DRAM[47433] = 8'b10110111;
DRAM[47434] = 8'b10110110;
DRAM[47435] = 8'b10111011;
DRAM[47436] = 8'b10111100;
DRAM[47437] = 8'b10110101;
DRAM[47438] = 8'b10101110;
DRAM[47439] = 8'b10101011;
DRAM[47440] = 8'b10101011;
DRAM[47441] = 8'b10100000;
DRAM[47442] = 8'b10010001;
DRAM[47443] = 8'b10000111;
DRAM[47444] = 8'b10001101;
DRAM[47445] = 8'b10011100;
DRAM[47446] = 8'b10100111;
DRAM[47447] = 8'b10101010;
DRAM[47448] = 8'b10010011;
DRAM[47449] = 8'b10010111;
DRAM[47450] = 8'b10010010;
DRAM[47451] = 8'b10001011;
DRAM[47452] = 8'b10001010;
DRAM[47453] = 8'b10000000;
DRAM[47454] = 8'b1111001;
DRAM[47455] = 8'b1111110;
DRAM[47456] = 8'b10000100;
DRAM[47457] = 8'b10001101;
DRAM[47458] = 8'b10000101;
DRAM[47459] = 8'b1110011;
DRAM[47460] = 8'b1111011;
DRAM[47461] = 8'b10010001;
DRAM[47462] = 8'b10001011;
DRAM[47463] = 8'b1110001;
DRAM[47464] = 8'b10000001;
DRAM[47465] = 8'b10001010;
DRAM[47466] = 8'b10010011;
DRAM[47467] = 8'b10011001;
DRAM[47468] = 8'b10011100;
DRAM[47469] = 8'b10011100;
DRAM[47470] = 8'b10010101;
DRAM[47471] = 8'b10001101;
DRAM[47472] = 8'b1110001;
DRAM[47473] = 8'b1101100;
DRAM[47474] = 8'b1111000;
DRAM[47475] = 8'b10010110;
DRAM[47476] = 8'b10101000;
DRAM[47477] = 8'b10100110;
DRAM[47478] = 8'b10100001;
DRAM[47479] = 8'b10100011;
DRAM[47480] = 8'b10011110;
DRAM[47481] = 8'b10011100;
DRAM[47482] = 8'b10001111;
DRAM[47483] = 8'b1111101;
DRAM[47484] = 8'b1110010;
DRAM[47485] = 8'b1110001;
DRAM[47486] = 8'b1101111;
DRAM[47487] = 8'b1101001;
DRAM[47488] = 8'b1100011;
DRAM[47489] = 8'b1010100;
DRAM[47490] = 8'b1000111;
DRAM[47491] = 8'b1000111;
DRAM[47492] = 8'b1001100;
DRAM[47493] = 8'b1001100;
DRAM[47494] = 8'b1000010;
DRAM[47495] = 8'b111000;
DRAM[47496] = 8'b110100;
DRAM[47497] = 8'b101010;
DRAM[47498] = 8'b100000;
DRAM[47499] = 8'b11110;
DRAM[47500] = 8'b11110;
DRAM[47501] = 8'b11001;
DRAM[47502] = 8'b1101;
DRAM[47503] = 8'b100;
DRAM[47504] = 8'b100;
DRAM[47505] = 8'b1;
DRAM[47506] = 8'b0;
DRAM[47507] = 8'b0;
DRAM[47508] = 8'b1;
DRAM[47509] = 8'b10;
DRAM[47510] = 8'b100;
DRAM[47511] = 8'b110;
DRAM[47512] = 8'b0;
DRAM[47513] = 8'b1;
DRAM[47514] = 8'b0;
DRAM[47515] = 8'b0;
DRAM[47516] = 8'b1010;
DRAM[47517] = 8'b1110;
DRAM[47518] = 8'b1100;
DRAM[47519] = 8'b10001;
DRAM[47520] = 8'b1011;
DRAM[47521] = 8'b11110;
DRAM[47522] = 8'b101011;
DRAM[47523] = 8'b110101;
DRAM[47524] = 8'b1000011;
DRAM[47525] = 8'b1001100;
DRAM[47526] = 8'b1010101;
DRAM[47527] = 8'b1100101;
DRAM[47528] = 8'b1101010;
DRAM[47529] = 8'b1110101;
DRAM[47530] = 8'b10000010;
DRAM[47531] = 8'b10001101;
DRAM[47532] = 8'b10011001;
DRAM[47533] = 8'b10101010;
DRAM[47534] = 8'b10111100;
DRAM[47535] = 8'b11001000;
DRAM[47536] = 8'b11000000;
DRAM[47537] = 8'b10111110;
DRAM[47538] = 8'b10111101;
DRAM[47539] = 8'b11000001;
DRAM[47540] = 8'b11001101;
DRAM[47541] = 8'b11011011;
DRAM[47542] = 8'b11100111;
DRAM[47543] = 8'b11101110;
DRAM[47544] = 8'b11110100;
DRAM[47545] = 8'b11110110;
DRAM[47546] = 8'b11111010;
DRAM[47547] = 8'b11111101;
DRAM[47548] = 8'b11111110;
DRAM[47549] = 8'b11111110;
DRAM[47550] = 8'b11111100;
DRAM[47551] = 8'b11111011;
DRAM[47552] = 8'b11111111;
DRAM[47553] = 8'b11111011;
DRAM[47554] = 8'b11110010;
DRAM[47555] = 8'b11101111;
DRAM[47556] = 8'b11101100;
DRAM[47557] = 8'b11100000;
DRAM[47558] = 8'b11001101;
DRAM[47559] = 8'b10111100;
DRAM[47560] = 8'b10110010;
DRAM[47561] = 8'b10100100;
DRAM[47562] = 8'b10011011;
DRAM[47563] = 8'b10011101;
DRAM[47564] = 8'b10011110;
DRAM[47565] = 8'b10011000;
DRAM[47566] = 8'b10010011;
DRAM[47567] = 8'b10010011;
DRAM[47568] = 8'b10001100;
DRAM[47569] = 8'b10001001;
DRAM[47570] = 8'b10000101;
DRAM[47571] = 8'b10000011;
DRAM[47572] = 8'b10000010;
DRAM[47573] = 8'b10000001;
DRAM[47574] = 8'b1111111;
DRAM[47575] = 8'b1111101;
DRAM[47576] = 8'b1111010;
DRAM[47577] = 8'b1111011;
DRAM[47578] = 8'b1111011;
DRAM[47579] = 8'b1111100;
DRAM[47580] = 8'b1111011;
DRAM[47581] = 8'b1111010;
DRAM[47582] = 8'b1111001;
DRAM[47583] = 8'b1111000;
DRAM[47584] = 8'b1111000;
DRAM[47585] = 8'b1111000;
DRAM[47586] = 8'b1111001;
DRAM[47587] = 8'b1111010;
DRAM[47588] = 8'b1111010;
DRAM[47589] = 8'b1111011;
DRAM[47590] = 8'b1111100;
DRAM[47591] = 8'b1111100;
DRAM[47592] = 8'b10000000;
DRAM[47593] = 8'b10000000;
DRAM[47594] = 8'b10000000;
DRAM[47595] = 8'b1111110;
DRAM[47596] = 8'b1111101;
DRAM[47597] = 8'b1111110;
DRAM[47598] = 8'b10000001;
DRAM[47599] = 8'b10000100;
DRAM[47600] = 8'b10000010;
DRAM[47601] = 8'b10000011;
DRAM[47602] = 8'b10000011;
DRAM[47603] = 8'b10000100;
DRAM[47604] = 8'b10000110;
DRAM[47605] = 8'b10001000;
DRAM[47606] = 8'b10001010;
DRAM[47607] = 8'b10001011;
DRAM[47608] = 8'b10001011;
DRAM[47609] = 8'b10001011;
DRAM[47610] = 8'b10001011;
DRAM[47611] = 8'b10001010;
DRAM[47612] = 8'b10001010;
DRAM[47613] = 8'b10001010;
DRAM[47614] = 8'b10001001;
DRAM[47615] = 8'b10001001;
DRAM[47616] = 8'b10001001;
DRAM[47617] = 8'b10001000;
DRAM[47618] = 8'b10000111;
DRAM[47619] = 8'b10001000;
DRAM[47620] = 8'b10001010;
DRAM[47621] = 8'b10001100;
DRAM[47622] = 8'b10001011;
DRAM[47623] = 8'b10001001;
DRAM[47624] = 8'b10001011;
DRAM[47625] = 8'b10001100;
DRAM[47626] = 8'b10001101;
DRAM[47627] = 8'b10001110;
DRAM[47628] = 8'b10001111;
DRAM[47629] = 8'b10010000;
DRAM[47630] = 8'b10010001;
DRAM[47631] = 8'b10010010;
DRAM[47632] = 8'b10010001;
DRAM[47633] = 8'b10010001;
DRAM[47634] = 8'b10010010;
DRAM[47635] = 8'b10010011;
DRAM[47636] = 8'b10010100;
DRAM[47637] = 8'b10010101;
DRAM[47638] = 8'b10010110;
DRAM[47639] = 8'b10010110;
DRAM[47640] = 8'b10010111;
DRAM[47641] = 8'b10011011;
DRAM[47642] = 8'b10011001;
DRAM[47643] = 8'b10011101;
DRAM[47644] = 8'b10100110;
DRAM[47645] = 8'b10101000;
DRAM[47646] = 8'b10101011;
DRAM[47647] = 8'b10111001;
DRAM[47648] = 8'b10111000;
DRAM[47649] = 8'b11001110;
DRAM[47650] = 8'b11101000;
DRAM[47651] = 8'b11111000;
DRAM[47652] = 8'b11111011;
DRAM[47653] = 8'b11111010;
DRAM[47654] = 8'b11111100;
DRAM[47655] = 8'b11111111;
DRAM[47656] = 8'b11111100;
DRAM[47657] = 8'b11111100;
DRAM[47658] = 8'b11111100;
DRAM[47659] = 8'b11111100;
DRAM[47660] = 8'b11111100;
DRAM[47661] = 8'b11111101;
DRAM[47662] = 8'b11111101;
DRAM[47663] = 8'b11111101;
DRAM[47664] = 8'b11111100;
DRAM[47665] = 8'b11111000;
DRAM[47666] = 8'b11110001;
DRAM[47667] = 8'b11101011;
DRAM[47668] = 8'b11100110;
DRAM[47669] = 8'b11100101;
DRAM[47670] = 8'b11100101;
DRAM[47671] = 8'b11100101;
DRAM[47672] = 8'b11100011;
DRAM[47673] = 8'b11100001;
DRAM[47674] = 8'b11011110;
DRAM[47675] = 8'b11011100;
DRAM[47676] = 8'b11011010;
DRAM[47677] = 8'b11011001;
DRAM[47678] = 8'b11011001;
DRAM[47679] = 8'b11011001;
DRAM[47680] = 8'b11001110;
DRAM[47681] = 8'b11010000;
DRAM[47682] = 8'b11010100;
DRAM[47683] = 8'b11010100;
DRAM[47684] = 8'b11001100;
DRAM[47685] = 8'b11000011;
DRAM[47686] = 8'b11000001;
DRAM[47687] = 8'b11000100;
DRAM[47688] = 8'b10111001;
DRAM[47689] = 8'b10110001;
DRAM[47690] = 8'b10101101;
DRAM[47691] = 8'b10110011;
DRAM[47692] = 8'b10111001;
DRAM[47693] = 8'b10110101;
DRAM[47694] = 8'b10101001;
DRAM[47695] = 8'b10100000;
DRAM[47696] = 8'b10011111;
DRAM[47697] = 8'b10010111;
DRAM[47698] = 8'b10010010;
DRAM[47699] = 8'b10010001;
DRAM[47700] = 8'b10010011;
DRAM[47701] = 8'b10010110;
DRAM[47702] = 8'b10011100;
DRAM[47703] = 8'b10100011;
DRAM[47704] = 8'b10010001;
DRAM[47705] = 8'b10011100;
DRAM[47706] = 8'b10011011;
DRAM[47707] = 8'b10010001;
DRAM[47708] = 8'b10001010;
DRAM[47709] = 8'b1111110;
DRAM[47710] = 8'b1111000;
DRAM[47711] = 8'b10000000;
DRAM[47712] = 8'b10001110;
DRAM[47713] = 8'b1111100;
DRAM[47714] = 8'b1110110;
DRAM[47715] = 8'b10000011;
DRAM[47716] = 8'b10001000;
DRAM[47717] = 8'b1111101;
DRAM[47718] = 8'b1111001;
DRAM[47719] = 8'b10000000;
DRAM[47720] = 8'b1110111;
DRAM[47721] = 8'b1111110;
DRAM[47722] = 8'b10001000;
DRAM[47723] = 8'b10010010;
DRAM[47724] = 8'b10011100;
DRAM[47725] = 8'b10100001;
DRAM[47726] = 8'b10011011;
DRAM[47727] = 8'b10010001;
DRAM[47728] = 8'b10000110;
DRAM[47729] = 8'b1111100;
DRAM[47730] = 8'b1111100;
DRAM[47731] = 8'b10001010;
DRAM[47732] = 8'b10010010;
DRAM[47733] = 8'b10010001;
DRAM[47734] = 8'b10010111;
DRAM[47735] = 8'b10100011;
DRAM[47736] = 8'b10011011;
DRAM[47737] = 8'b10010010;
DRAM[47738] = 8'b10001001;
DRAM[47739] = 8'b10000001;
DRAM[47740] = 8'b1110110;
DRAM[47741] = 8'b1101010;
DRAM[47742] = 8'b1100100;
DRAM[47743] = 8'b1100100;
DRAM[47744] = 8'b1011000;
DRAM[47745] = 8'b1000101;
DRAM[47746] = 8'b111001;
DRAM[47747] = 8'b1000001;
DRAM[47748] = 8'b1001011;
DRAM[47749] = 8'b1001000;
DRAM[47750] = 8'b111100;
DRAM[47751] = 8'b110100;
DRAM[47752] = 8'b101000;
DRAM[47753] = 8'b11101;
DRAM[47754] = 8'b10001;
DRAM[47755] = 8'b1100;
DRAM[47756] = 8'b1101;
DRAM[47757] = 8'b1011;
DRAM[47758] = 8'b10;
DRAM[47759] = 8'b0;
DRAM[47760] = 8'b10;
DRAM[47761] = 8'b0;
DRAM[47762] = 8'b0;
DRAM[47763] = 8'b101;
DRAM[47764] = 8'b101;
DRAM[47765] = 8'b0;
DRAM[47766] = 8'b0;
DRAM[47767] = 8'b10;
DRAM[47768] = 8'b0;
DRAM[47769] = 8'b1100;
DRAM[47770] = 8'b1001;
DRAM[47771] = 8'b1;
DRAM[47772] = 8'b1100;
DRAM[47773] = 8'b11010;
DRAM[47774] = 8'b11101;
DRAM[47775] = 8'b11110;
DRAM[47776] = 8'b10010;
DRAM[47777] = 8'b101010;
DRAM[47778] = 8'b111100;
DRAM[47779] = 8'b1000110;
DRAM[47780] = 8'b1001111;
DRAM[47781] = 8'b1010011;
DRAM[47782] = 8'b1011110;
DRAM[47783] = 8'b1110010;
DRAM[47784] = 8'b1110101;
DRAM[47785] = 8'b10000011;
DRAM[47786] = 8'b10010000;
DRAM[47787] = 8'b10010111;
DRAM[47788] = 8'b10100011;
DRAM[47789] = 8'b10110100;
DRAM[47790] = 8'b11000001;
DRAM[47791] = 8'b11000101;
DRAM[47792] = 8'b10110011;
DRAM[47793] = 8'b10110011;
DRAM[47794] = 8'b10111000;
DRAM[47795] = 8'b11000100;
DRAM[47796] = 8'b11010110;
DRAM[47797] = 8'b11100110;
DRAM[47798] = 8'b11101111;
DRAM[47799] = 8'b11110011;
DRAM[47800] = 8'b11110110;
DRAM[47801] = 8'b11111000;
DRAM[47802] = 8'b11111011;
DRAM[47803] = 8'b11111110;
DRAM[47804] = 8'b11111110;
DRAM[47805] = 8'b11111110;
DRAM[47806] = 8'b11111101;
DRAM[47807] = 8'b11111011;
DRAM[47808] = 8'b11111111;
DRAM[47809] = 8'b11111101;
DRAM[47810] = 8'b11110111;
DRAM[47811] = 8'b11110101;
DRAM[47812] = 8'b11110010;
DRAM[47813] = 8'b11100100;
DRAM[47814] = 8'b11001101;
DRAM[47815] = 8'b10111010;
DRAM[47816] = 8'b10110011;
DRAM[47817] = 8'b10100101;
DRAM[47818] = 8'b10010111;
DRAM[47819] = 8'b10010011;
DRAM[47820] = 8'b10011000;
DRAM[47821] = 8'b10011011;
DRAM[47822] = 8'b10010111;
DRAM[47823] = 8'b10010001;
DRAM[47824] = 8'b10001010;
DRAM[47825] = 8'b10000111;
DRAM[47826] = 8'b10000100;
DRAM[47827] = 8'b10000010;
DRAM[47828] = 8'b10000001;
DRAM[47829] = 8'b1111111;
DRAM[47830] = 8'b1111101;
DRAM[47831] = 8'b1111011;
DRAM[47832] = 8'b1111000;
DRAM[47833] = 8'b1111000;
DRAM[47834] = 8'b1111001;
DRAM[47835] = 8'b1111001;
DRAM[47836] = 8'b1111000;
DRAM[47837] = 8'b1111000;
DRAM[47838] = 8'b1110111;
DRAM[47839] = 8'b1110110;
DRAM[47840] = 8'b1111000;
DRAM[47841] = 8'b1111000;
DRAM[47842] = 8'b1111001;
DRAM[47843] = 8'b1111010;
DRAM[47844] = 8'b1111010;
DRAM[47845] = 8'b1111011;
DRAM[47846] = 8'b1111100;
DRAM[47847] = 8'b1111100;
DRAM[47848] = 8'b1111110;
DRAM[47849] = 8'b1111111;
DRAM[47850] = 8'b10000000;
DRAM[47851] = 8'b1111111;
DRAM[47852] = 8'b1111110;
DRAM[47853] = 8'b1111111;
DRAM[47854] = 8'b10000001;
DRAM[47855] = 8'b10000011;
DRAM[47856] = 8'b10000010;
DRAM[47857] = 8'b10000011;
DRAM[47858] = 8'b10000011;
DRAM[47859] = 8'b10000100;
DRAM[47860] = 8'b10000110;
DRAM[47861] = 8'b10000111;
DRAM[47862] = 8'b10001001;
DRAM[47863] = 8'b10001010;
DRAM[47864] = 8'b10001100;
DRAM[47865] = 8'b10001100;
DRAM[47866] = 8'b10001011;
DRAM[47867] = 8'b10001011;
DRAM[47868] = 8'b10001010;
DRAM[47869] = 8'b10001010;
DRAM[47870] = 8'b10001010;
DRAM[47871] = 8'b10001010;
DRAM[47872] = 8'b10001010;
DRAM[47873] = 8'b10001001;
DRAM[47874] = 8'b10001001;
DRAM[47875] = 8'b10001010;
DRAM[47876] = 8'b10001100;
DRAM[47877] = 8'b10001101;
DRAM[47878] = 8'b10001101;
DRAM[47879] = 8'b10001100;
DRAM[47880] = 8'b10001010;
DRAM[47881] = 8'b10001011;
DRAM[47882] = 8'b10001100;
DRAM[47883] = 8'b10001101;
DRAM[47884] = 8'b10001110;
DRAM[47885] = 8'b10001111;
DRAM[47886] = 8'b10010000;
DRAM[47887] = 8'b10010001;
DRAM[47888] = 8'b10010000;
DRAM[47889] = 8'b10010000;
DRAM[47890] = 8'b10010001;
DRAM[47891] = 8'b10010010;
DRAM[47892] = 8'b10010011;
DRAM[47893] = 8'b10010100;
DRAM[47894] = 8'b10010101;
DRAM[47895] = 8'b10010110;
DRAM[47896] = 8'b10010100;
DRAM[47897] = 8'b10011001;
DRAM[47898] = 8'b10011001;
DRAM[47899] = 8'b10011101;
DRAM[47900] = 8'b10100111;
DRAM[47901] = 8'b10101001;
DRAM[47902] = 8'b10101110;
DRAM[47903] = 8'b10111101;
DRAM[47904] = 8'b11001100;
DRAM[47905] = 8'b11100001;
DRAM[47906] = 8'b11111000;
DRAM[47907] = 8'b11111111;
DRAM[47908] = 8'b11111111;
DRAM[47909] = 8'b11111101;
DRAM[47910] = 8'b11111110;
DRAM[47911] = 8'b11111111;
DRAM[47912] = 8'b11111100;
DRAM[47913] = 8'b11111101;
DRAM[47914] = 8'b11111101;
DRAM[47915] = 8'b11111101;
DRAM[47916] = 8'b11111101;
DRAM[47917] = 8'b11111101;
DRAM[47918] = 8'b11111101;
DRAM[47919] = 8'b11111100;
DRAM[47920] = 8'b11111010;
DRAM[47921] = 8'b11110101;
DRAM[47922] = 8'b11101110;
DRAM[47923] = 8'b11101000;
DRAM[47924] = 8'b11100100;
DRAM[47925] = 8'b11100011;
DRAM[47926] = 8'b11100010;
DRAM[47927] = 8'b11100010;
DRAM[47928] = 8'b11100010;
DRAM[47929] = 8'b11100000;
DRAM[47930] = 8'b11011110;
DRAM[47931] = 8'b11011101;
DRAM[47932] = 8'b11011101;
DRAM[47933] = 8'b11011110;
DRAM[47934] = 8'b11011110;
DRAM[47935] = 8'b11011110;
DRAM[47936] = 8'b11010010;
DRAM[47937] = 8'b11011001;
DRAM[47938] = 8'b11011111;
DRAM[47939] = 8'b11011110;
DRAM[47940] = 8'b11010011;
DRAM[47941] = 8'b11000111;
DRAM[47942] = 8'b11000001;
DRAM[47943] = 8'b11000001;
DRAM[47944] = 8'b10111000;
DRAM[47945] = 8'b10110001;
DRAM[47946] = 8'b10101100;
DRAM[47947] = 8'b10101111;
DRAM[47948] = 8'b10110100;
DRAM[47949] = 8'b10110001;
DRAM[47950] = 8'b10100111;
DRAM[47951] = 8'b10011101;
DRAM[47952] = 8'b10011001;
DRAM[47953] = 8'b10010001;
DRAM[47954] = 8'b10001111;
DRAM[47955] = 8'b10010101;
DRAM[47956] = 8'b10010110;
DRAM[47957] = 8'b10010001;
DRAM[47958] = 8'b10010001;
DRAM[47959] = 8'b10010111;
DRAM[47960] = 8'b10010101;
DRAM[47961] = 8'b10100011;
DRAM[47962] = 8'b10100010;
DRAM[47963] = 8'b10011000;
DRAM[47964] = 8'b10010011;
DRAM[47965] = 8'b10001010;
DRAM[47966] = 8'b10000100;
DRAM[47967] = 8'b10001001;
DRAM[47968] = 8'b10000000;
DRAM[47969] = 8'b1110000;
DRAM[47970] = 8'b1110110;
DRAM[47971] = 8'b10001011;
DRAM[47972] = 8'b10000110;
DRAM[47973] = 8'b1101110;
DRAM[47974] = 8'b1110101;
DRAM[47975] = 8'b10010011;
DRAM[47976] = 8'b1110011;
DRAM[47977] = 8'b1111010;
DRAM[47978] = 8'b10000010;
DRAM[47979] = 8'b10001010;
DRAM[47980] = 8'b10010100;
DRAM[47981] = 8'b10011100;
DRAM[47982] = 8'b10011100;
DRAM[47983] = 8'b10010110;
DRAM[47984] = 8'b10011001;
DRAM[47985] = 8'b10001100;
DRAM[47986] = 8'b10000000;
DRAM[47987] = 8'b1111100;
DRAM[47988] = 8'b1111010;
DRAM[47989] = 8'b1111100;
DRAM[47990] = 8'b10001101;
DRAM[47991] = 8'b10100001;
DRAM[47992] = 8'b10010100;
DRAM[47993] = 8'b10010010;
DRAM[47994] = 8'b10001111;
DRAM[47995] = 8'b10001001;
DRAM[47996] = 8'b1111101;
DRAM[47997] = 8'b1101101;
DRAM[47998] = 8'b1011111;
DRAM[47999] = 8'b1011000;
DRAM[48000] = 8'b1001110;
DRAM[48001] = 8'b1000000;
DRAM[48002] = 8'b111011;
DRAM[48003] = 8'b1000111;
DRAM[48004] = 8'b1001110;
DRAM[48005] = 8'b1000010;
DRAM[48006] = 8'b110001;
DRAM[48007] = 8'b101000;
DRAM[48008] = 8'b10101;
DRAM[48009] = 8'b10001;
DRAM[48010] = 8'b1001;
DRAM[48011] = 8'b11;
DRAM[48012] = 8'b11;
DRAM[48013] = 8'b111;
DRAM[48014] = 8'b111;
DRAM[48015] = 8'b100;
DRAM[48016] = 8'b111;
DRAM[48017] = 8'b10;
DRAM[48018] = 8'b100;
DRAM[48019] = 8'b1101;
DRAM[48020] = 8'b1100;
DRAM[48021] = 8'b11;
DRAM[48022] = 8'b11;
DRAM[48023] = 8'b1010;
DRAM[48024] = 8'b10111;
DRAM[48025] = 8'b100000;
DRAM[48026] = 8'b11011;
DRAM[48027] = 8'b10101;
DRAM[48028] = 8'b100010;
DRAM[48029] = 8'b110000;
DRAM[48030] = 8'b110111;
DRAM[48031] = 8'b111111;
DRAM[48032] = 8'b111001;
DRAM[48033] = 8'b1001011;
DRAM[48034] = 8'b1010111;
DRAM[48035] = 8'b1011101;
DRAM[48036] = 8'b1100010;
DRAM[48037] = 8'b1100001;
DRAM[48038] = 8'b1101001;
DRAM[48039] = 8'b1111101;
DRAM[48040] = 8'b10000001;
DRAM[48041] = 8'b10010110;
DRAM[48042] = 8'b10100111;
DRAM[48043] = 8'b10101010;
DRAM[48044] = 8'b10101100;
DRAM[48045] = 8'b10110010;
DRAM[48046] = 8'b10110100;
DRAM[48047] = 8'b10110000;
DRAM[48048] = 8'b10101101;
DRAM[48049] = 8'b10110010;
DRAM[48050] = 8'b10111100;
DRAM[48051] = 8'b11001010;
DRAM[48052] = 8'b11011001;
DRAM[48053] = 8'b11100101;
DRAM[48054] = 8'b11101101;
DRAM[48055] = 8'b11110001;
DRAM[48056] = 8'b11111001;
DRAM[48057] = 8'b11111010;
DRAM[48058] = 8'b11111100;
DRAM[48059] = 8'b11111110;
DRAM[48060] = 8'b11111110;
DRAM[48061] = 8'b11111110;
DRAM[48062] = 8'b11111101;
DRAM[48063] = 8'b11111100;
DRAM[48064] = 8'b11111100;
DRAM[48065] = 8'b11111110;
DRAM[48066] = 8'b11111101;
DRAM[48067] = 8'b11110100;
DRAM[48068] = 8'b11100100;
DRAM[48069] = 8'b11010001;
DRAM[48070] = 8'b11000010;
DRAM[48071] = 8'b10111010;
DRAM[48072] = 8'b10110011;
DRAM[48073] = 8'b10101010;
DRAM[48074] = 8'b10011100;
DRAM[48075] = 8'b10010010;
DRAM[48076] = 8'b10010100;
DRAM[48077] = 8'b10011001;
DRAM[48078] = 8'b10010110;
DRAM[48079] = 8'b10001110;
DRAM[48080] = 8'b10001000;
DRAM[48081] = 8'b10000101;
DRAM[48082] = 8'b10000010;
DRAM[48083] = 8'b10000000;
DRAM[48084] = 8'b1111111;
DRAM[48085] = 8'b1111110;
DRAM[48086] = 8'b1111011;
DRAM[48087] = 8'b1111001;
DRAM[48088] = 8'b1110110;
DRAM[48089] = 8'b1110110;
DRAM[48090] = 8'b1110111;
DRAM[48091] = 8'b1110111;
DRAM[48092] = 8'b1110111;
DRAM[48093] = 8'b1110110;
DRAM[48094] = 8'b1110110;
DRAM[48095] = 8'b1110110;
DRAM[48096] = 8'b1111000;
DRAM[48097] = 8'b1111000;
DRAM[48098] = 8'b1111001;
DRAM[48099] = 8'b1111010;
DRAM[48100] = 8'b1111010;
DRAM[48101] = 8'b1111011;
DRAM[48102] = 8'b1111100;
DRAM[48103] = 8'b1111100;
DRAM[48104] = 8'b1111100;
DRAM[48105] = 8'b1111110;
DRAM[48106] = 8'b10000000;
DRAM[48107] = 8'b10000000;
DRAM[48108] = 8'b1111111;
DRAM[48109] = 8'b1111111;
DRAM[48110] = 8'b10000000;
DRAM[48111] = 8'b10000010;
DRAM[48112] = 8'b10000011;
DRAM[48113] = 8'b10000011;
DRAM[48114] = 8'b10000011;
DRAM[48115] = 8'b10000100;
DRAM[48116] = 8'b10000101;
DRAM[48117] = 8'b10000111;
DRAM[48118] = 8'b10001000;
DRAM[48119] = 8'b10001001;
DRAM[48120] = 8'b10001100;
DRAM[48121] = 8'b10001011;
DRAM[48122] = 8'b10001011;
DRAM[48123] = 8'b10001011;
DRAM[48124] = 8'b10001010;
DRAM[48125] = 8'b10001010;
DRAM[48126] = 8'b10001010;
DRAM[48127] = 8'b10001010;
DRAM[48128] = 8'b10001010;
DRAM[48129] = 8'b10001001;
DRAM[48130] = 8'b10001000;
DRAM[48131] = 8'b10001010;
DRAM[48132] = 8'b10001100;
DRAM[48133] = 8'b10001110;
DRAM[48134] = 8'b10001101;
DRAM[48135] = 8'b10001100;
DRAM[48136] = 8'b10001011;
DRAM[48137] = 8'b10001011;
DRAM[48138] = 8'b10001100;
DRAM[48139] = 8'b10001101;
DRAM[48140] = 8'b10001111;
DRAM[48141] = 8'b10010000;
DRAM[48142] = 8'b10010001;
DRAM[48143] = 8'b10010001;
DRAM[48144] = 8'b10010001;
DRAM[48145] = 8'b10010001;
DRAM[48146] = 8'b10010010;
DRAM[48147] = 8'b10010010;
DRAM[48148] = 8'b10010011;
DRAM[48149] = 8'b10010100;
DRAM[48150] = 8'b10010101;
DRAM[48151] = 8'b10010101;
DRAM[48152] = 8'b10010100;
DRAM[48153] = 8'b10011001;
DRAM[48154] = 8'b10011000;
DRAM[48155] = 8'b10011010;
DRAM[48156] = 8'b10100011;
DRAM[48157] = 8'b10100101;
DRAM[48158] = 8'b10101100;
DRAM[48159] = 8'b10111101;
DRAM[48160] = 8'b11011111;
DRAM[48161] = 8'b11101111;
DRAM[48162] = 8'b11111110;
DRAM[48163] = 8'b11111111;
DRAM[48164] = 8'b11111110;
DRAM[48165] = 8'b11111111;
DRAM[48166] = 8'b11111111;
DRAM[48167] = 8'b11111110;
DRAM[48168] = 8'b11111101;
DRAM[48169] = 8'b11111110;
DRAM[48170] = 8'b11111110;
DRAM[48171] = 8'b11111111;
DRAM[48172] = 8'b11111110;
DRAM[48173] = 8'b11111101;
DRAM[48174] = 8'b11111100;
DRAM[48175] = 8'b11111011;
DRAM[48176] = 8'b11111010;
DRAM[48177] = 8'b11110110;
DRAM[48178] = 8'b11110001;
DRAM[48179] = 8'b11101110;
DRAM[48180] = 8'b11101100;
DRAM[48181] = 8'b11101011;
DRAM[48182] = 8'b11101000;
DRAM[48183] = 8'b11100101;
DRAM[48184] = 8'b11011110;
DRAM[48185] = 8'b11011011;
DRAM[48186] = 8'b11011001;
DRAM[48187] = 8'b11011001;
DRAM[48188] = 8'b11011011;
DRAM[48189] = 8'b11011101;
DRAM[48190] = 8'b11011101;
DRAM[48191] = 8'b11011100;
DRAM[48192] = 8'b11011100;
DRAM[48193] = 8'b11011111;
DRAM[48194] = 8'b11100000;
DRAM[48195] = 8'b11011010;
DRAM[48196] = 8'b11010001;
DRAM[48197] = 8'b11001010;
DRAM[48198] = 8'b11001000;
DRAM[48199] = 8'b11001000;
DRAM[48200] = 8'b10111010;
DRAM[48201] = 8'b10110111;
DRAM[48202] = 8'b10110011;
DRAM[48203] = 8'b10101111;
DRAM[48204] = 8'b10101100;
DRAM[48205] = 8'b10101010;
DRAM[48206] = 8'b10100101;
DRAM[48207] = 8'b10100001;
DRAM[48208] = 8'b10011111;
DRAM[48209] = 8'b10001110;
DRAM[48210] = 8'b10000010;
DRAM[48211] = 8'b10000101;
DRAM[48212] = 8'b10001010;
DRAM[48213] = 8'b10001100;
DRAM[48214] = 8'b10010001;
DRAM[48215] = 8'b10011001;
DRAM[48216] = 8'b10001101;
DRAM[48217] = 8'b10011000;
DRAM[48218] = 8'b10010101;
DRAM[48219] = 8'b10001111;
DRAM[48220] = 8'b10010011;
DRAM[48221] = 8'b10010001;
DRAM[48222] = 8'b10001000;
DRAM[48223] = 8'b10000111;
DRAM[48224] = 8'b1110111;
DRAM[48225] = 8'b10000101;
DRAM[48226] = 8'b10001000;
DRAM[48227] = 8'b1111001;
DRAM[48228] = 8'b1110000;
DRAM[48229] = 8'b1110110;
DRAM[48230] = 8'b1111010;
DRAM[48231] = 8'b1110111;
DRAM[48232] = 8'b1110000;
DRAM[48233] = 8'b1111000;
DRAM[48234] = 8'b1111111;
DRAM[48235] = 8'b10000010;
DRAM[48236] = 8'b10001000;
DRAM[48237] = 8'b10010010;
DRAM[48238] = 8'b10011001;
DRAM[48239] = 8'b10011100;
DRAM[48240] = 8'b10010110;
DRAM[48241] = 8'b10001101;
DRAM[48242] = 8'b10000011;
DRAM[48243] = 8'b1111011;
DRAM[48244] = 8'b1110010;
DRAM[48245] = 8'b1110001;
DRAM[48246] = 8'b10000000;
DRAM[48247] = 8'b10010010;
DRAM[48248] = 8'b10001101;
DRAM[48249] = 8'b10010101;
DRAM[48250] = 8'b10010011;
DRAM[48251] = 8'b10000111;
DRAM[48252] = 8'b1111101;
DRAM[48253] = 8'b1111000;
DRAM[48254] = 8'b1101100;
DRAM[48255] = 8'b1011101;
DRAM[48256] = 8'b1010100;
DRAM[48257] = 8'b1001011;
DRAM[48258] = 8'b1001010;
DRAM[48259] = 8'b1010000;
DRAM[48260] = 8'b1001101;
DRAM[48261] = 8'b111110;
DRAM[48262] = 8'b101110;
DRAM[48263] = 8'b101000;
DRAM[48264] = 8'b10110;
DRAM[48265] = 8'b11001;
DRAM[48266] = 8'b10101;
DRAM[48267] = 8'b1100;
DRAM[48268] = 8'b1000;
DRAM[48269] = 8'b1101;
DRAM[48270] = 8'b10010;
DRAM[48271] = 8'b10011;
DRAM[48272] = 8'b1110;
DRAM[48273] = 8'b1011;
DRAM[48274] = 8'b10000;
DRAM[48275] = 8'b11000;
DRAM[48276] = 8'b11010;
DRAM[48277] = 8'b10111;
DRAM[48278] = 8'b11011;
DRAM[48279] = 8'b100101;
DRAM[48280] = 8'b101001;
DRAM[48281] = 8'b101011;
DRAM[48282] = 8'b101011;
DRAM[48283] = 8'b110100;
DRAM[48284] = 8'b1000010;
DRAM[48285] = 8'b1000011;
DRAM[48286] = 8'b1000110;
DRAM[48287] = 8'b1010100;
DRAM[48288] = 8'b1011001;
DRAM[48289] = 8'b1100001;
DRAM[48290] = 8'b1100100;
DRAM[48291] = 8'b1101001;
DRAM[48292] = 8'b1110010;
DRAM[48293] = 8'b1110010;
DRAM[48294] = 8'b1111000;
DRAM[48295] = 8'b10001010;
DRAM[48296] = 8'b10011001;
DRAM[48297] = 8'b10101100;
DRAM[48298] = 8'b10111010;
DRAM[48299] = 8'b10110100;
DRAM[48300] = 8'b10101001;
DRAM[48301] = 8'b10100101;
DRAM[48302] = 8'b10100011;
DRAM[48303] = 8'b10100000;
DRAM[48304] = 8'b10100110;
DRAM[48305] = 8'b10110000;
DRAM[48306] = 8'b10111110;
DRAM[48307] = 8'b11001010;
DRAM[48308] = 8'b11010010;
DRAM[48309] = 8'b11011011;
DRAM[48310] = 8'b11100101;
DRAM[48311] = 8'b11101101;
DRAM[48312] = 8'b11111001;
DRAM[48313] = 8'b11111010;
DRAM[48314] = 8'b11111100;
DRAM[48315] = 8'b11111101;
DRAM[48316] = 8'b11111110;
DRAM[48317] = 8'b11111110;
DRAM[48318] = 8'b11111101;
DRAM[48319] = 8'b11111100;
DRAM[48320] = 8'b11111100;
DRAM[48321] = 8'b11111110;
DRAM[48322] = 8'b11111110;
DRAM[48323] = 8'b11110101;
DRAM[48324] = 8'b11100011;
DRAM[48325] = 8'b11001110;
DRAM[48326] = 8'b10111100;
DRAM[48327] = 8'b10110011;
DRAM[48328] = 8'b10101100;
DRAM[48329] = 8'b10101000;
DRAM[48330] = 8'b10011111;
DRAM[48331] = 8'b10010100;
DRAM[48332] = 8'b10010001;
DRAM[48333] = 8'b10010011;
DRAM[48334] = 8'b10010001;
DRAM[48335] = 8'b10001100;
DRAM[48336] = 8'b10000110;
DRAM[48337] = 8'b10000011;
DRAM[48338] = 8'b10000000;
DRAM[48339] = 8'b1111110;
DRAM[48340] = 8'b1111101;
DRAM[48341] = 8'b1111011;
DRAM[48342] = 8'b1111001;
DRAM[48343] = 8'b1110111;
DRAM[48344] = 8'b1110110;
DRAM[48345] = 8'b1110110;
DRAM[48346] = 8'b1110101;
DRAM[48347] = 8'b1110101;
DRAM[48348] = 8'b1110101;
DRAM[48349] = 8'b1110110;
DRAM[48350] = 8'b1110110;
DRAM[48351] = 8'b1110110;
DRAM[48352] = 8'b1111000;
DRAM[48353] = 8'b1111000;
DRAM[48354] = 8'b1111001;
DRAM[48355] = 8'b1111010;
DRAM[48356] = 8'b1111010;
DRAM[48357] = 8'b1111011;
DRAM[48358] = 8'b1111100;
DRAM[48359] = 8'b1111100;
DRAM[48360] = 8'b1111011;
DRAM[48361] = 8'b1111101;
DRAM[48362] = 8'b1111111;
DRAM[48363] = 8'b1111111;
DRAM[48364] = 8'b1111111;
DRAM[48365] = 8'b1111111;
DRAM[48366] = 8'b10000000;
DRAM[48367] = 8'b10000010;
DRAM[48368] = 8'b10000011;
DRAM[48369] = 8'b10000011;
DRAM[48370] = 8'b10000011;
DRAM[48371] = 8'b10000011;
DRAM[48372] = 8'b10000101;
DRAM[48373] = 8'b10000110;
DRAM[48374] = 8'b10001000;
DRAM[48375] = 8'b10001000;
DRAM[48376] = 8'b10001011;
DRAM[48377] = 8'b10001011;
DRAM[48378] = 8'b10001010;
DRAM[48379] = 8'b10001010;
DRAM[48380] = 8'b10001010;
DRAM[48381] = 8'b10001001;
DRAM[48382] = 8'b10001001;
DRAM[48383] = 8'b10001001;
DRAM[48384] = 8'b10001000;
DRAM[48385] = 8'b10000111;
DRAM[48386] = 8'b10000110;
DRAM[48387] = 8'b10001000;
DRAM[48388] = 8'b10001011;
DRAM[48389] = 8'b10001100;
DRAM[48390] = 8'b10001100;
DRAM[48391] = 8'b10001011;
DRAM[48392] = 8'b10001101;
DRAM[48393] = 8'b10001101;
DRAM[48394] = 8'b10001110;
DRAM[48395] = 8'b10001111;
DRAM[48396] = 8'b10010000;
DRAM[48397] = 8'b10010001;
DRAM[48398] = 8'b10010010;
DRAM[48399] = 8'b10010011;
DRAM[48400] = 8'b10010011;
DRAM[48401] = 8'b10010011;
DRAM[48402] = 8'b10010011;
DRAM[48403] = 8'b10010011;
DRAM[48404] = 8'b10010100;
DRAM[48405] = 8'b10010100;
DRAM[48406] = 8'b10010100;
DRAM[48407] = 8'b10010100;
DRAM[48408] = 8'b10010110;
DRAM[48409] = 8'b10011001;
DRAM[48410] = 8'b10010110;
DRAM[48411] = 8'b10010101;
DRAM[48412] = 8'b10011100;
DRAM[48413] = 8'b10011111;
DRAM[48414] = 8'b10101010;
DRAM[48415] = 8'b10111110;
DRAM[48416] = 8'b11100110;
DRAM[48417] = 8'b11110010;
DRAM[48418] = 8'b11111011;
DRAM[48419] = 8'b11111010;
DRAM[48420] = 8'b11111001;
DRAM[48421] = 8'b11111110;
DRAM[48422] = 8'b11111111;
DRAM[48423] = 8'b11111011;
DRAM[48424] = 8'b11111110;
DRAM[48425] = 8'b11111110;
DRAM[48426] = 8'b11111111;
DRAM[48427] = 8'b11111111;
DRAM[48428] = 8'b11111110;
DRAM[48429] = 8'b11111011;
DRAM[48430] = 8'b11111001;
DRAM[48431] = 8'b11111000;
DRAM[48432] = 8'b11110011;
DRAM[48433] = 8'b11110000;
DRAM[48434] = 8'b11101101;
DRAM[48435] = 8'b11101100;
DRAM[48436] = 8'b11101101;
DRAM[48437] = 8'b11101011;
DRAM[48438] = 8'b11100110;
DRAM[48439] = 8'b11100001;
DRAM[48440] = 8'b11011101;
DRAM[48441] = 8'b11011001;
DRAM[48442] = 8'b11010110;
DRAM[48443] = 8'b11010111;
DRAM[48444] = 8'b11011011;
DRAM[48445] = 8'b11011110;
DRAM[48446] = 8'b11011101;
DRAM[48447] = 8'b11011100;
DRAM[48448] = 8'b11011111;
DRAM[48449] = 8'b11011101;
DRAM[48450] = 8'b11010111;
DRAM[48451] = 8'b11001101;
DRAM[48452] = 8'b11001000;
DRAM[48453] = 8'b11001011;
DRAM[48454] = 8'b11001111;
DRAM[48455] = 8'b11010000;
DRAM[48456] = 8'b10111100;
DRAM[48457] = 8'b10111110;
DRAM[48458] = 8'b10111010;
DRAM[48459] = 8'b10101111;
DRAM[48460] = 8'b10100110;
DRAM[48461] = 8'b10100011;
DRAM[48462] = 8'b10100010;
DRAM[48463] = 8'b10100000;
DRAM[48464] = 8'b10010010;
DRAM[48465] = 8'b10001000;
DRAM[48466] = 8'b10000001;
DRAM[48467] = 8'b10000100;
DRAM[48468] = 8'b10001010;
DRAM[48469] = 8'b10001101;
DRAM[48470] = 8'b10001101;
DRAM[48471] = 8'b10001101;
DRAM[48472] = 8'b10000001;
DRAM[48473] = 8'b10001010;
DRAM[48474] = 8'b10000101;
DRAM[48475] = 8'b10000010;
DRAM[48476] = 8'b10001101;
DRAM[48477] = 8'b10010010;
DRAM[48478] = 8'b10001010;
DRAM[48479] = 8'b10000101;
DRAM[48480] = 8'b10001001;
DRAM[48481] = 8'b10000110;
DRAM[48482] = 8'b1111100;
DRAM[48483] = 8'b1110010;
DRAM[48484] = 8'b1110010;
DRAM[48485] = 8'b1111000;
DRAM[48486] = 8'b1110010;
DRAM[48487] = 8'b1100110;
DRAM[48488] = 8'b1101111;
DRAM[48489] = 8'b1110110;
DRAM[48490] = 8'b1111010;
DRAM[48491] = 8'b1111001;
DRAM[48492] = 8'b1111100;
DRAM[48493] = 8'b10000111;
DRAM[48494] = 8'b10010011;
DRAM[48495] = 8'b10011001;
DRAM[48496] = 8'b10001111;
DRAM[48497] = 8'b10001111;
DRAM[48498] = 8'b10001111;
DRAM[48499] = 8'b10001000;
DRAM[48500] = 8'b1111000;
DRAM[48501] = 8'b1101010;
DRAM[48502] = 8'b1101010;
DRAM[48503] = 8'b1110001;
DRAM[48504] = 8'b10001000;
DRAM[48505] = 8'b10010001;
DRAM[48506] = 8'b10001111;
DRAM[48507] = 8'b10000011;
DRAM[48508] = 8'b1111110;
DRAM[48509] = 8'b10000010;
DRAM[48510] = 8'b1111101;
DRAM[48511] = 8'b1110001;
DRAM[48512] = 8'b1100101;
DRAM[48513] = 8'b1100001;
DRAM[48514] = 8'b1011011;
DRAM[48515] = 8'b1010101;
DRAM[48516] = 8'b1001111;
DRAM[48517] = 8'b1000111;
DRAM[48518] = 8'b111110;
DRAM[48519] = 8'b111000;
DRAM[48520] = 8'b100100;
DRAM[48521] = 8'b101011;
DRAM[48522] = 8'b101011;
DRAM[48523] = 8'b100010;
DRAM[48524] = 8'b11111;
DRAM[48525] = 8'b100110;
DRAM[48526] = 8'b101101;
DRAM[48527] = 8'b101101;
DRAM[48528] = 8'b100100;
DRAM[48529] = 8'b100111;
DRAM[48530] = 8'b101001;
DRAM[48531] = 8'b101010;
DRAM[48532] = 8'b101001;
DRAM[48533] = 8'b101011;
DRAM[48534] = 8'b110001;
DRAM[48535] = 8'b110110;
DRAM[48536] = 8'b110011;
DRAM[48537] = 8'b110110;
DRAM[48538] = 8'b111101;
DRAM[48539] = 8'b1001110;
DRAM[48540] = 8'b1011100;
DRAM[48541] = 8'b1010100;
DRAM[48542] = 8'b1010000;
DRAM[48543] = 8'b1011101;
DRAM[48544] = 8'b1101010;
DRAM[48545] = 8'b1101010;
DRAM[48546] = 8'b1101001;
DRAM[48547] = 8'b1110010;
DRAM[48548] = 8'b10000011;
DRAM[48549] = 8'b10001000;
DRAM[48550] = 8'b10010001;
DRAM[48551] = 8'b10100100;
DRAM[48552] = 8'b10110111;
DRAM[48553] = 8'b10111010;
DRAM[48554] = 8'b10111000;
DRAM[48555] = 8'b10101101;
DRAM[48556] = 8'b10011110;
DRAM[48557] = 8'b10010111;
DRAM[48558] = 8'b10011100;
DRAM[48559] = 8'b10100011;
DRAM[48560] = 8'b10100110;
DRAM[48561] = 8'b10110010;
DRAM[48562] = 8'b11000001;
DRAM[48563] = 8'b11001011;
DRAM[48564] = 8'b11010000;
DRAM[48565] = 8'b11011001;
DRAM[48566] = 8'b11100111;
DRAM[48567] = 8'b11110010;
DRAM[48568] = 8'b11111000;
DRAM[48569] = 8'b11111001;
DRAM[48570] = 8'b11111010;
DRAM[48571] = 8'b11111100;
DRAM[48572] = 8'b11111101;
DRAM[48573] = 8'b11111101;
DRAM[48574] = 8'b11111101;
DRAM[48575] = 8'b11111101;
DRAM[48576] = 8'b11111111;
DRAM[48577] = 8'b11111101;
DRAM[48578] = 8'b11111011;
DRAM[48579] = 8'b11111011;
DRAM[48580] = 8'b11110101;
DRAM[48581] = 8'b11100010;
DRAM[48582] = 8'b11000100;
DRAM[48583] = 8'b10101101;
DRAM[48584] = 8'b10100100;
DRAM[48585] = 8'b10011111;
DRAM[48586] = 8'b10011001;
DRAM[48587] = 8'b10010011;
DRAM[48588] = 8'b10001111;
DRAM[48589] = 8'b10001101;
DRAM[48590] = 8'b10001100;
DRAM[48591] = 8'b10001011;
DRAM[48592] = 8'b10000100;
DRAM[48593] = 8'b10000001;
DRAM[48594] = 8'b1111110;
DRAM[48595] = 8'b1111100;
DRAM[48596] = 8'b1111011;
DRAM[48597] = 8'b1111010;
DRAM[48598] = 8'b1110111;
DRAM[48599] = 8'b1110101;
DRAM[48600] = 8'b1110100;
DRAM[48601] = 8'b1110100;
DRAM[48602] = 8'b1110011;
DRAM[48603] = 8'b1110011;
DRAM[48604] = 8'b1110100;
DRAM[48605] = 8'b1110100;
DRAM[48606] = 8'b1110101;
DRAM[48607] = 8'b1110110;
DRAM[48608] = 8'b1111000;
DRAM[48609] = 8'b1111000;
DRAM[48610] = 8'b1111001;
DRAM[48611] = 8'b1111010;
DRAM[48612] = 8'b1111010;
DRAM[48613] = 8'b1111011;
DRAM[48614] = 8'b1111100;
DRAM[48615] = 8'b1111100;
DRAM[48616] = 8'b1111011;
DRAM[48617] = 8'b1111101;
DRAM[48618] = 8'b1111110;
DRAM[48619] = 8'b1111110;
DRAM[48620] = 8'b1111101;
DRAM[48621] = 8'b1111110;
DRAM[48622] = 8'b10000001;
DRAM[48623] = 8'b10000011;
DRAM[48624] = 8'b10000011;
DRAM[48625] = 8'b10000011;
DRAM[48626] = 8'b10000011;
DRAM[48627] = 8'b10000011;
DRAM[48628] = 8'b10000100;
DRAM[48629] = 8'b10000101;
DRAM[48630] = 8'b10000111;
DRAM[48631] = 8'b10001000;
DRAM[48632] = 8'b10001001;
DRAM[48633] = 8'b10001001;
DRAM[48634] = 8'b10001001;
DRAM[48635] = 8'b10001000;
DRAM[48636] = 8'b10001000;
DRAM[48637] = 8'b10001000;
DRAM[48638] = 8'b10000111;
DRAM[48639] = 8'b10000111;
DRAM[48640] = 8'b10001000;
DRAM[48641] = 8'b10000111;
DRAM[48642] = 8'b10000111;
DRAM[48643] = 8'b10001001;
DRAM[48644] = 8'b10001100;
DRAM[48645] = 8'b10001110;
DRAM[48646] = 8'b10001101;
DRAM[48647] = 8'b10001100;
DRAM[48648] = 8'b10001111;
DRAM[48649] = 8'b10001111;
DRAM[48650] = 8'b10010000;
DRAM[48651] = 8'b10010001;
DRAM[48652] = 8'b10010010;
DRAM[48653] = 8'b10010100;
DRAM[48654] = 8'b10010100;
DRAM[48655] = 8'b10010101;
DRAM[48656] = 8'b10010101;
DRAM[48657] = 8'b10010101;
DRAM[48658] = 8'b10010101;
DRAM[48659] = 8'b10010101;
DRAM[48660] = 8'b10010100;
DRAM[48661] = 8'b10010100;
DRAM[48662] = 8'b10010100;
DRAM[48663] = 8'b10010100;
DRAM[48664] = 8'b10010101;
DRAM[48665] = 8'b10011000;
DRAM[48666] = 8'b10010011;
DRAM[48667] = 8'b10010010;
DRAM[48668] = 8'b10011010;
DRAM[48669] = 8'b10100010;
DRAM[48670] = 8'b10110010;
DRAM[48671] = 8'b11001010;
DRAM[48672] = 8'b11101000;
DRAM[48673] = 8'b11110110;
DRAM[48674] = 8'b11111110;
DRAM[48675] = 8'b11111010;
DRAM[48676] = 8'b11111000;
DRAM[48677] = 8'b11111100;
DRAM[48678] = 8'b11111110;
DRAM[48679] = 8'b11111011;
DRAM[48680] = 8'b11111101;
DRAM[48681] = 8'b11111110;
DRAM[48682] = 8'b11111110;
DRAM[48683] = 8'b11111101;
DRAM[48684] = 8'b11111011;
DRAM[48685] = 8'b11111000;
DRAM[48686] = 8'b11110101;
DRAM[48687] = 8'b11110011;
DRAM[48688] = 8'b11101101;
DRAM[48689] = 8'b11101001;
DRAM[48690] = 8'b11100100;
DRAM[48691] = 8'b11100011;
DRAM[48692] = 8'b11100100;
DRAM[48693] = 8'b11100011;
DRAM[48694] = 8'b11011110;
DRAM[48695] = 8'b11011001;
DRAM[48696] = 8'b11011101;
DRAM[48697] = 8'b11011001;
DRAM[48698] = 8'b11010101;
DRAM[48699] = 8'b11010110;
DRAM[48700] = 8'b11011011;
DRAM[48701] = 8'b11011110;
DRAM[48702] = 8'b11011110;
DRAM[48703] = 8'b11011011;
DRAM[48704] = 8'b11011000;
DRAM[48705] = 8'b11011000;
DRAM[48706] = 8'b11010010;
DRAM[48707] = 8'b11001011;
DRAM[48708] = 8'b11001010;
DRAM[48709] = 8'b11001110;
DRAM[48710] = 8'b11001101;
DRAM[48711] = 8'b11000111;
DRAM[48712] = 8'b10111101;
DRAM[48713] = 8'b11000001;
DRAM[48714] = 8'b10111100;
DRAM[48715] = 8'b10110000;
DRAM[48716] = 8'b10100100;
DRAM[48717] = 8'b10011111;
DRAM[48718] = 8'b10011100;
DRAM[48719] = 8'b10010111;
DRAM[48720] = 8'b10000101;
DRAM[48721] = 8'b10001001;
DRAM[48722] = 8'b10001010;
DRAM[48723] = 8'b10001010;
DRAM[48724] = 8'b10001010;
DRAM[48725] = 8'b10001001;
DRAM[48726] = 8'b10000011;
DRAM[48727] = 8'b1111011;
DRAM[48728] = 8'b1111010;
DRAM[48729] = 8'b10000100;
DRAM[48730] = 8'b10000000;
DRAM[48731] = 8'b1111101;
DRAM[48732] = 8'b10001011;
DRAM[48733] = 8'b10010100;
DRAM[48734] = 8'b10001111;
DRAM[48735] = 8'b10001010;
DRAM[48736] = 8'b10010100;
DRAM[48737] = 8'b1111010;
DRAM[48738] = 8'b1101101;
DRAM[48739] = 8'b1110111;
DRAM[48740] = 8'b1111010;
DRAM[48741] = 8'b1101101;
DRAM[48742] = 8'b1100111;
DRAM[48743] = 8'b1101110;
DRAM[48744] = 8'b1110100;
DRAM[48745] = 8'b1110110;
DRAM[48746] = 8'b1110101;
DRAM[48747] = 8'b1110010;
DRAM[48748] = 8'b1110101;
DRAM[48749] = 8'b1111110;
DRAM[48750] = 8'b10000101;
DRAM[48751] = 8'b10000111;
DRAM[48752] = 8'b10001100;
DRAM[48753] = 8'b10010010;
DRAM[48754] = 8'b10010111;
DRAM[48755] = 8'b10010011;
DRAM[48756] = 8'b10000010;
DRAM[48757] = 8'b1101111;
DRAM[48758] = 8'b1100110;
DRAM[48759] = 8'b1100110;
DRAM[48760] = 8'b10000000;
DRAM[48761] = 8'b10000100;
DRAM[48762] = 8'b10001001;
DRAM[48763] = 8'b10001011;
DRAM[48764] = 8'b10001010;
DRAM[48765] = 8'b10000111;
DRAM[48766] = 8'b10000001;
DRAM[48767] = 8'b1111100;
DRAM[48768] = 8'b1110001;
DRAM[48769] = 8'b1110001;
DRAM[48770] = 8'b1101010;
DRAM[48771] = 8'b1100000;
DRAM[48772] = 8'b1011110;
DRAM[48773] = 8'b1100000;
DRAM[48774] = 8'b1011000;
DRAM[48775] = 8'b1001010;
DRAM[48776] = 8'b111011;
DRAM[48777] = 8'b1000001;
DRAM[48778] = 8'b1000000;
DRAM[48779] = 8'b111011;
DRAM[48780] = 8'b111110;
DRAM[48781] = 8'b1001000;
DRAM[48782] = 8'b1001010;
DRAM[48783] = 8'b1000100;
DRAM[48784] = 8'b111001;
DRAM[48785] = 8'b1000011;
DRAM[48786] = 8'b1000101;
DRAM[48787] = 8'b111100;
DRAM[48788] = 8'b111001;
DRAM[48789] = 8'b111110;
DRAM[48790] = 8'b1000001;
DRAM[48791] = 8'b111111;
DRAM[48792] = 8'b111111;
DRAM[48793] = 8'b1000111;
DRAM[48794] = 8'b1001010;
DRAM[48795] = 8'b1010010;
DRAM[48796] = 8'b1011111;
DRAM[48797] = 8'b1100000;
DRAM[48798] = 8'b1011110;
DRAM[48799] = 8'b1100111;
DRAM[48800] = 8'b1110011;
DRAM[48801] = 8'b1110011;
DRAM[48802] = 8'b1110011;
DRAM[48803] = 8'b10000000;
DRAM[48804] = 8'b10010011;
DRAM[48805] = 8'b10011010;
DRAM[48806] = 8'b10100110;
DRAM[48807] = 8'b10111011;
DRAM[48808] = 8'b11000100;
DRAM[48809] = 8'b10110100;
DRAM[48810] = 8'b10100101;
DRAM[48811] = 8'b10011101;
DRAM[48812] = 8'b10010101;
DRAM[48813] = 8'b10010010;
DRAM[48814] = 8'b10011100;
DRAM[48815] = 8'b10101011;
DRAM[48816] = 8'b10101111;
DRAM[48817] = 8'b10110110;
DRAM[48818] = 8'b11000000;
DRAM[48819] = 8'b11001001;
DRAM[48820] = 8'b11010001;
DRAM[48821] = 8'b11011101;
DRAM[48822] = 8'b11101100;
DRAM[48823] = 8'b11110110;
DRAM[48824] = 8'b11110110;
DRAM[48825] = 8'b11110111;
DRAM[48826] = 8'b11111001;
DRAM[48827] = 8'b11111010;
DRAM[48828] = 8'b11111100;
DRAM[48829] = 8'b11111101;
DRAM[48830] = 8'b11111110;
DRAM[48831] = 8'b11111110;
DRAM[48832] = 8'b11111111;
DRAM[48833] = 8'b11111100;
DRAM[48834] = 8'b11111011;
DRAM[48835] = 8'b11111101;
DRAM[48836] = 8'b11111100;
DRAM[48837] = 8'b11101101;
DRAM[48838] = 8'b11010011;
DRAM[48839] = 8'b10111111;
DRAM[48840] = 8'b10101010;
DRAM[48841] = 8'b10011100;
DRAM[48842] = 8'b10010010;
DRAM[48843] = 8'b10010010;
DRAM[48844] = 8'b10010000;
DRAM[48845] = 8'b10001010;
DRAM[48846] = 8'b10000111;
DRAM[48847] = 8'b10001001;
DRAM[48848] = 8'b10000011;
DRAM[48849] = 8'b10000000;
DRAM[48850] = 8'b1111100;
DRAM[48851] = 8'b1111010;
DRAM[48852] = 8'b1111001;
DRAM[48853] = 8'b1111000;
DRAM[48854] = 8'b1110110;
DRAM[48855] = 8'b1110100;
DRAM[48856] = 8'b1110010;
DRAM[48857] = 8'b1110001;
DRAM[48858] = 8'b1110001;
DRAM[48859] = 8'b1110000;
DRAM[48860] = 8'b1110001;
DRAM[48861] = 8'b1110010;
DRAM[48862] = 8'b1110011;
DRAM[48863] = 8'b1110100;
DRAM[48864] = 8'b1111000;
DRAM[48865] = 8'b1111000;
DRAM[48866] = 8'b1111001;
DRAM[48867] = 8'b1111010;
DRAM[48868] = 8'b1111010;
DRAM[48869] = 8'b1111011;
DRAM[48870] = 8'b1111100;
DRAM[48871] = 8'b1111100;
DRAM[48872] = 8'b1111100;
DRAM[48873] = 8'b1111101;
DRAM[48874] = 8'b1111101;
DRAM[48875] = 8'b1111100;
DRAM[48876] = 8'b1111100;
DRAM[48877] = 8'b1111110;
DRAM[48878] = 8'b10000010;
DRAM[48879] = 8'b10000101;
DRAM[48880] = 8'b10000011;
DRAM[48881] = 8'b10000011;
DRAM[48882] = 8'b10000011;
DRAM[48883] = 8'b10000011;
DRAM[48884] = 8'b10000100;
DRAM[48885] = 8'b10000101;
DRAM[48886] = 8'b10000110;
DRAM[48887] = 8'b10000111;
DRAM[48888] = 8'b10001000;
DRAM[48889] = 8'b10001000;
DRAM[48890] = 8'b10000111;
DRAM[48891] = 8'b10000111;
DRAM[48892] = 8'b10000111;
DRAM[48893] = 8'b10000110;
DRAM[48894] = 8'b10000110;
DRAM[48895] = 8'b10000110;
DRAM[48896] = 8'b10001011;
DRAM[48897] = 8'b10001010;
DRAM[48898] = 8'b10001010;
DRAM[48899] = 8'b10001100;
DRAM[48900] = 8'b10001111;
DRAM[48901] = 8'b10010001;
DRAM[48902] = 8'b10010001;
DRAM[48903] = 8'b10010000;
DRAM[48904] = 8'b10010000;
DRAM[48905] = 8'b10010001;
DRAM[48906] = 8'b10010010;
DRAM[48907] = 8'b10010011;
DRAM[48908] = 8'b10010100;
DRAM[48909] = 8'b10010101;
DRAM[48910] = 8'b10010110;
DRAM[48911] = 8'b10010110;
DRAM[48912] = 8'b10010111;
DRAM[48913] = 8'b10010111;
DRAM[48914] = 8'b10010110;
DRAM[48915] = 8'b10010110;
DRAM[48916] = 8'b10010101;
DRAM[48917] = 8'b10010100;
DRAM[48918] = 8'b10010011;
DRAM[48919] = 8'b10010011;
DRAM[48920] = 8'b10010011;
DRAM[48921] = 8'b10010110;
DRAM[48922] = 8'b10010001;
DRAM[48923] = 8'b10010001;
DRAM[48924] = 8'b10011101;
DRAM[48925] = 8'b10101001;
DRAM[48926] = 8'b10111110;
DRAM[48927] = 8'b11011010;
DRAM[48928] = 8'b11101100;
DRAM[48929] = 8'b11111110;
DRAM[48930] = 8'b11111111;
DRAM[48931] = 8'b11111111;
DRAM[48932] = 8'b11111010;
DRAM[48933] = 8'b11111100;
DRAM[48934] = 8'b11111111;
DRAM[48935] = 8'b11111100;
DRAM[48936] = 8'b11111100;
DRAM[48937] = 8'b11111100;
DRAM[48938] = 8'b11111100;
DRAM[48939] = 8'b11111011;
DRAM[48940] = 8'b11111001;
DRAM[48941] = 8'b11110101;
DRAM[48942] = 8'b11110001;
DRAM[48943] = 8'b11101111;
DRAM[48944] = 8'b11101111;
DRAM[48945] = 8'b11101001;
DRAM[48946] = 8'b11100010;
DRAM[48947] = 8'b11100000;
DRAM[48948] = 8'b11100001;
DRAM[48949] = 8'b11100000;
DRAM[48950] = 8'b11011100;
DRAM[48951] = 8'b11010111;
DRAM[48952] = 8'b11011010;
DRAM[48953] = 8'b11010101;
DRAM[48954] = 8'b11010001;
DRAM[48955] = 8'b11010011;
DRAM[48956] = 8'b11011000;
DRAM[48957] = 8'b11011011;
DRAM[48958] = 8'b11011010;
DRAM[48959] = 8'b11010111;
DRAM[48960] = 8'b11010000;
DRAM[48961] = 8'b11010100;
DRAM[48962] = 8'b11010110;
DRAM[48963] = 8'b11010100;
DRAM[48964] = 8'b11010101;
DRAM[48965] = 8'b11010010;
DRAM[48966] = 8'b11000101;
DRAM[48967] = 8'b10110110;
DRAM[48968] = 8'b10111101;
DRAM[48969] = 8'b11000000;
DRAM[48970] = 8'b10111100;
DRAM[48971] = 8'b10101111;
DRAM[48972] = 8'b10100101;
DRAM[48973] = 8'b10011111;
DRAM[48974] = 8'b10010111;
DRAM[48975] = 8'b10001110;
DRAM[48976] = 8'b10010000;
DRAM[48977] = 8'b10010101;
DRAM[48978] = 8'b10010000;
DRAM[48979] = 8'b10000001;
DRAM[48980] = 8'b1111001;
DRAM[48981] = 8'b1111100;
DRAM[48982] = 8'b1111111;
DRAM[48983] = 8'b1111100;
DRAM[48984] = 8'b1110111;
DRAM[48985] = 8'b10000100;
DRAM[48986] = 8'b10000001;
DRAM[48987] = 8'b1111100;
DRAM[48988] = 8'b10001001;
DRAM[48989] = 8'b10010100;
DRAM[48990] = 8'b10010001;
DRAM[48991] = 8'b10001111;
DRAM[48992] = 8'b10001001;
DRAM[48993] = 8'b10000110;
DRAM[48994] = 8'b1111101;
DRAM[48995] = 8'b1110001;
DRAM[48996] = 8'b1101010;
DRAM[48997] = 8'b1101010;
DRAM[48998] = 8'b1101010;
DRAM[48999] = 8'b1101010;
DRAM[49000] = 8'b1111011;
DRAM[49001] = 8'b1111000;
DRAM[49002] = 8'b1110011;
DRAM[49003] = 8'b1101111;
DRAM[49004] = 8'b1110010;
DRAM[49005] = 8'b1111000;
DRAM[49006] = 8'b1111000;
DRAM[49007] = 8'b1110011;
DRAM[49008] = 8'b10000100;
DRAM[49009] = 8'b10001100;
DRAM[49010] = 8'b10010100;
DRAM[49011] = 8'b10010100;
DRAM[49012] = 8'b10001001;
DRAM[49013] = 8'b1111101;
DRAM[49014] = 8'b1111001;
DRAM[49015] = 8'b1111011;
DRAM[49016] = 8'b1111000;
DRAM[49017] = 8'b1111001;
DRAM[49018] = 8'b10000111;
DRAM[49019] = 8'b10011001;
DRAM[49020] = 8'b10011001;
DRAM[49021] = 8'b10000111;
DRAM[49022] = 8'b1111001;
DRAM[49023] = 8'b1111001;
DRAM[49024] = 8'b1110001;
DRAM[49025] = 8'b1110111;
DRAM[49026] = 8'b1110011;
DRAM[49027] = 8'b1101100;
DRAM[49028] = 8'b1110001;
DRAM[49029] = 8'b1111000;
DRAM[49030] = 8'b1101010;
DRAM[49031] = 8'b1010010;
DRAM[49032] = 8'b1010111;
DRAM[49033] = 8'b1010111;
DRAM[49034] = 8'b1010010;
DRAM[49035] = 8'b1001100;
DRAM[49036] = 8'b1010010;
DRAM[49037] = 8'b1011011;
DRAM[49038] = 8'b1010110;
DRAM[49039] = 8'b1000111;
DRAM[49040] = 8'b111010;
DRAM[49041] = 8'b1001011;
DRAM[49042] = 8'b1010000;
DRAM[49043] = 8'b1000111;
DRAM[49044] = 8'b1000101;
DRAM[49045] = 8'b1001111;
DRAM[49046] = 8'b1010011;
DRAM[49047] = 8'b1001100;
DRAM[49048] = 8'b1001001;
DRAM[49049] = 8'b1010011;
DRAM[49050] = 8'b1001101;
DRAM[49051] = 8'b1000100;
DRAM[49052] = 8'b1010000;
DRAM[49053] = 8'b1100001;
DRAM[49054] = 8'b1101001;
DRAM[49055] = 8'b1101111;
DRAM[49056] = 8'b1111001;
DRAM[49057] = 8'b1111010;
DRAM[49058] = 8'b1111100;
DRAM[49059] = 8'b10001001;
DRAM[49060] = 8'b10011010;
DRAM[49061] = 8'b10011111;
DRAM[49062] = 8'b10101011;
DRAM[49063] = 8'b11000011;
DRAM[49064] = 8'b11000001;
DRAM[49065] = 8'b10100110;
DRAM[49066] = 8'b10010010;
DRAM[49067] = 8'b10010010;
DRAM[49068] = 8'b10010100;
DRAM[49069] = 8'b10010010;
DRAM[49070] = 8'b10011100;
DRAM[49071] = 8'b10101100;
DRAM[49072] = 8'b10110011;
DRAM[49073] = 8'b10110101;
DRAM[49074] = 8'b10111010;
DRAM[49075] = 8'b11000010;
DRAM[49076] = 8'b11001101;
DRAM[49077] = 8'b11011011;
DRAM[49078] = 8'b11101001;
DRAM[49079] = 8'b11110001;
DRAM[49080] = 8'b11110101;
DRAM[49081] = 8'b11110110;
DRAM[49082] = 8'b11110111;
DRAM[49083] = 8'b11111001;
DRAM[49084] = 8'b11111011;
DRAM[49085] = 8'b11111101;
DRAM[49086] = 8'b11111110;
DRAM[49087] = 8'b11111111;
DRAM[49088] = 8'b11111000;
DRAM[49089] = 8'b11111011;
DRAM[49090] = 8'b11111110;
DRAM[49091] = 8'b11111011;
DRAM[49092] = 8'b11110010;
DRAM[49093] = 8'b11100110;
DRAM[49094] = 8'b11011101;
DRAM[49095] = 8'b11011001;
DRAM[49096] = 8'b10110111;
DRAM[49097] = 8'b10100000;
DRAM[49098] = 8'b10010000;
DRAM[49099] = 8'b10010010;
DRAM[49100] = 8'b10010011;
DRAM[49101] = 8'b10001001;
DRAM[49102] = 8'b10000011;
DRAM[49103] = 8'b10000110;
DRAM[49104] = 8'b10000010;
DRAM[49105] = 8'b1111111;
DRAM[49106] = 8'b1111100;
DRAM[49107] = 8'b1111001;
DRAM[49108] = 8'b1111001;
DRAM[49109] = 8'b1110111;
DRAM[49110] = 8'b1110101;
DRAM[49111] = 8'b1110011;
DRAM[49112] = 8'b1110000;
DRAM[49113] = 8'b1101111;
DRAM[49114] = 8'b1101110;
DRAM[49115] = 8'b1101110;
DRAM[49116] = 8'b1101110;
DRAM[49117] = 8'b1110000;
DRAM[49118] = 8'b1110010;
DRAM[49119] = 8'b1110011;
DRAM[49120] = 8'b1111000;
DRAM[49121] = 8'b1111000;
DRAM[49122] = 8'b1111001;
DRAM[49123] = 8'b1111010;
DRAM[49124] = 8'b1111010;
DRAM[49125] = 8'b1111011;
DRAM[49126] = 8'b1111100;
DRAM[49127] = 8'b1111100;
DRAM[49128] = 8'b1111101;
DRAM[49129] = 8'b1111101;
DRAM[49130] = 8'b1111100;
DRAM[49131] = 8'b1111011;
DRAM[49132] = 8'b1111011;
DRAM[49133] = 8'b1111101;
DRAM[49134] = 8'b10000010;
DRAM[49135] = 8'b10000110;
DRAM[49136] = 8'b10000011;
DRAM[49137] = 8'b10000011;
DRAM[49138] = 8'b10000011;
DRAM[49139] = 8'b10000011;
DRAM[49140] = 8'b10000011;
DRAM[49141] = 8'b10000101;
DRAM[49142] = 8'b10000110;
DRAM[49143] = 8'b10000110;
DRAM[49144] = 8'b10000111;
DRAM[49145] = 8'b10000111;
DRAM[49146] = 8'b10000110;
DRAM[49147] = 8'b10000110;
DRAM[49148] = 8'b10000110;
DRAM[49149] = 8'b10000101;
DRAM[49150] = 8'b10000101;
DRAM[49151] = 8'b10000101;
DRAM[49152] = 8'b10000111;
DRAM[49153] = 8'b10001000;
DRAM[49154] = 8'b10001001;
DRAM[49155] = 8'b10001011;
DRAM[49156] = 8'b10001101;
DRAM[49157] = 8'b10001110;
DRAM[49158] = 8'b10010000;
DRAM[49159] = 8'b10010000;
DRAM[49160] = 8'b10010101;
DRAM[49161] = 8'b10010010;
DRAM[49162] = 8'b10010001;
DRAM[49163] = 8'b10010001;
DRAM[49164] = 8'b10010011;
DRAM[49165] = 8'b10010110;
DRAM[49166] = 8'b10010111;
DRAM[49167] = 8'b10010110;
DRAM[49168] = 8'b10011001;
DRAM[49169] = 8'b10011001;
DRAM[49170] = 8'b10011000;
DRAM[49171] = 8'b10010110;
DRAM[49172] = 8'b10010110;
DRAM[49173] = 8'b10010110;
DRAM[49174] = 8'b10010110;
DRAM[49175] = 8'b10010110;
DRAM[49176] = 8'b10010001;
DRAM[49177] = 8'b10010110;
DRAM[49178] = 8'b10011111;
DRAM[49179] = 8'b10100010;
DRAM[49180] = 8'b10011110;
DRAM[49181] = 8'b10100100;
DRAM[49182] = 8'b11000111;
DRAM[49183] = 8'b11101101;
DRAM[49184] = 8'b11111100;
DRAM[49185] = 8'b11111100;
DRAM[49186] = 8'b11111110;
DRAM[49187] = 8'b11111111;
DRAM[49188] = 8'b11111111;
DRAM[49189] = 8'b11111111;
DRAM[49190] = 8'b11111111;
DRAM[49191] = 8'b11111111;
DRAM[49192] = 8'b11111111;
DRAM[49193] = 8'b11111101;
DRAM[49194] = 8'b11111011;
DRAM[49195] = 8'b11111000;
DRAM[49196] = 8'b11110101;
DRAM[49197] = 8'b11110100;
DRAM[49198] = 8'b11110100;
DRAM[49199] = 8'b11110011;
DRAM[49200] = 8'b11110000;
DRAM[49201] = 8'b11101110;
DRAM[49202] = 8'b11100011;
DRAM[49203] = 8'b11011101;
DRAM[49204] = 8'b11011111;
DRAM[49205] = 8'b11011010;
DRAM[49206] = 8'b11010111;
DRAM[49207] = 8'b11100001;
DRAM[49208] = 8'b11011010;
DRAM[49209] = 8'b11011100;
DRAM[49210] = 8'b11011111;
DRAM[49211] = 8'b11100000;
DRAM[49212] = 8'b11011111;
DRAM[49213] = 8'b11011100;
DRAM[49214] = 8'b11011000;
DRAM[49215] = 8'b11010110;
DRAM[49216] = 8'b11011000;
DRAM[49217] = 8'b11010010;
DRAM[49218] = 8'b11001101;
DRAM[49219] = 8'b11001011;
DRAM[49220] = 8'b11001100;
DRAM[49221] = 8'b11001100;
DRAM[49222] = 8'b11000111;
DRAM[49223] = 8'b11000011;
DRAM[49224] = 8'b10111010;
DRAM[49225] = 8'b10101011;
DRAM[49226] = 8'b10100010;
DRAM[49227] = 8'b10100100;
DRAM[49228] = 8'b10100111;
DRAM[49229] = 8'b10100001;
DRAM[49230] = 8'b10011001;
DRAM[49231] = 8'b10010100;
DRAM[49232] = 8'b10011101;
DRAM[49233] = 8'b10000110;
DRAM[49234] = 8'b1111011;
DRAM[49235] = 8'b10000101;
DRAM[49236] = 8'b10000110;
DRAM[49237] = 8'b1111000;
DRAM[49238] = 8'b1110011;
DRAM[49239] = 8'b1111100;
DRAM[49240] = 8'b1111110;
DRAM[49241] = 8'b1111101;
DRAM[49242] = 8'b1111101;
DRAM[49243] = 8'b10001101;
DRAM[49244] = 8'b10011110;
DRAM[49245] = 8'b10011001;
DRAM[49246] = 8'b10001111;
DRAM[49247] = 8'b10010001;
DRAM[49248] = 8'b10001000;
DRAM[49249] = 8'b10000100;
DRAM[49250] = 8'b1110111;
DRAM[49251] = 8'b1111100;
DRAM[49252] = 8'b1110011;
DRAM[49253] = 8'b1100010;
DRAM[49254] = 8'b1110011;
DRAM[49255] = 8'b10000000;
DRAM[49256] = 8'b1111111;
DRAM[49257] = 8'b1110111;
DRAM[49258] = 8'b1101100;
DRAM[49259] = 8'b1101000;
DRAM[49260] = 8'b1110000;
DRAM[49261] = 8'b1111001;
DRAM[49262] = 8'b1110101;
DRAM[49263] = 8'b1101011;
DRAM[49264] = 8'b1110110;
DRAM[49265] = 8'b1111101;
DRAM[49266] = 8'b10000110;
DRAM[49267] = 8'b10001000;
DRAM[49268] = 8'b10000110;
DRAM[49269] = 8'b10000011;
DRAM[49270] = 8'b10000011;
DRAM[49271] = 8'b10000110;
DRAM[49272] = 8'b1111011;
DRAM[49273] = 8'b1111100;
DRAM[49274] = 8'b10000010;
DRAM[49275] = 8'b10001101;
DRAM[49276] = 8'b10010101;
DRAM[49277] = 8'b10010101;
DRAM[49278] = 8'b10001100;
DRAM[49279] = 8'b10000011;
DRAM[49280] = 8'b1111011;
DRAM[49281] = 8'b10000000;
DRAM[49282] = 8'b10000001;
DRAM[49283] = 8'b1111011;
DRAM[49284] = 8'b1110101;
DRAM[49285] = 8'b1110011;
DRAM[49286] = 8'b1110000;
DRAM[49287] = 8'b1101101;
DRAM[49288] = 8'b1101011;
DRAM[49289] = 8'b1101011;
DRAM[49290] = 8'b1101000;
DRAM[49291] = 8'b1100011;
DRAM[49292] = 8'b1100001;
DRAM[49293] = 8'b1011110;
DRAM[49294] = 8'b1010110;
DRAM[49295] = 8'b1001101;
DRAM[49296] = 8'b1000111;
DRAM[49297] = 8'b1001110;
DRAM[49298] = 8'b1010100;
DRAM[49299] = 8'b1010010;
DRAM[49300] = 8'b1010000;
DRAM[49301] = 8'b1010011;
DRAM[49302] = 8'b1011011;
DRAM[49303] = 8'b1100001;
DRAM[49304] = 8'b1010100;
DRAM[49305] = 8'b1001101;
DRAM[49306] = 8'b1001110;
DRAM[49307] = 8'b1010001;
DRAM[49308] = 8'b1010010;
DRAM[49309] = 8'b1100010;
DRAM[49310] = 8'b1110010;
DRAM[49311] = 8'b1110010;
DRAM[49312] = 8'b10000010;
DRAM[49313] = 8'b1111011;
DRAM[49314] = 8'b10001100;
DRAM[49315] = 8'b10001110;
DRAM[49316] = 8'b10100100;
DRAM[49317] = 8'b10110010;
DRAM[49318] = 8'b10011101;
DRAM[49319] = 8'b10101001;
DRAM[49320] = 8'b10100111;
DRAM[49321] = 8'b10011101;
DRAM[49322] = 8'b10010110;
DRAM[49323] = 8'b10011000;
DRAM[49324] = 8'b10011100;
DRAM[49325] = 8'b10011110;
DRAM[49326] = 8'b10100000;
DRAM[49327] = 8'b10100010;
DRAM[49328] = 8'b10101001;
DRAM[49329] = 8'b10110100;
DRAM[49330] = 8'b11000011;
DRAM[49331] = 8'b11001101;
DRAM[49332] = 8'b11010100;
DRAM[49333] = 8'b11011101;
DRAM[49334] = 8'b11101011;
DRAM[49335] = 8'b11110110;
DRAM[49336] = 8'b11110110;
DRAM[49337] = 8'b11110111;
DRAM[49338] = 8'b11110111;
DRAM[49339] = 8'b11110111;
DRAM[49340] = 8'b11110111;
DRAM[49341] = 8'b11111001;
DRAM[49342] = 8'b11111101;
DRAM[49343] = 8'b11111111;
DRAM[49344] = 8'b11110110;
DRAM[49345] = 8'b11111011;
DRAM[49346] = 8'b11111010;
DRAM[49347] = 8'b11110100;
DRAM[49348] = 8'b11110010;
DRAM[49349] = 8'b11101111;
DRAM[49350] = 8'b11011111;
DRAM[49351] = 8'b11001100;
DRAM[49352] = 8'b10111010;
DRAM[49353] = 8'b10101111;
DRAM[49354] = 8'b10100011;
DRAM[49355] = 8'b10011011;
DRAM[49356] = 8'b10010011;
DRAM[49357] = 8'b10001001;
DRAM[49358] = 8'b10000101;
DRAM[49359] = 8'b10000101;
DRAM[49360] = 8'b1111111;
DRAM[49361] = 8'b1111110;
DRAM[49362] = 8'b1111101;
DRAM[49363] = 8'b1111010;
DRAM[49364] = 8'b1111000;
DRAM[49365] = 8'b1110110;
DRAM[49366] = 8'b1110100;
DRAM[49367] = 8'b1110011;
DRAM[49368] = 8'b1110001;
DRAM[49369] = 8'b1110000;
DRAM[49370] = 8'b1101111;
DRAM[49371] = 8'b1101111;
DRAM[49372] = 8'b1110000;
DRAM[49373] = 8'b1110010;
DRAM[49374] = 8'b1110011;
DRAM[49375] = 8'b1110101;
DRAM[49376] = 8'b1110100;
DRAM[49377] = 8'b1110101;
DRAM[49378] = 8'b1110111;
DRAM[49379] = 8'b1111000;
DRAM[49380] = 8'b1111001;
DRAM[49381] = 8'b1111010;
DRAM[49382] = 8'b1111010;
DRAM[49383] = 8'b1111010;
DRAM[49384] = 8'b1111010;
DRAM[49385] = 8'b1111010;
DRAM[49386] = 8'b1111011;
DRAM[49387] = 8'b1111100;
DRAM[49388] = 8'b1111101;
DRAM[49389] = 8'b1111111;
DRAM[49390] = 8'b10000000;
DRAM[49391] = 8'b10000001;
DRAM[49392] = 8'b10000011;
DRAM[49393] = 8'b10000011;
DRAM[49394] = 8'b10000011;
DRAM[49395] = 8'b10000100;
DRAM[49396] = 8'b10000100;
DRAM[49397] = 8'b10000101;
DRAM[49398] = 8'b10000101;
DRAM[49399] = 8'b10000110;
DRAM[49400] = 8'b10000100;
DRAM[49401] = 8'b10000100;
DRAM[49402] = 8'b10000100;
DRAM[49403] = 8'b10000101;
DRAM[49404] = 8'b10000110;
DRAM[49405] = 8'b10000110;
DRAM[49406] = 8'b10000110;
DRAM[49407] = 8'b10000111;
DRAM[49408] = 8'b10001001;
DRAM[49409] = 8'b10001010;
DRAM[49410] = 8'b10001011;
DRAM[49411] = 8'b10001101;
DRAM[49412] = 8'b10001111;
DRAM[49413] = 8'b10010000;
DRAM[49414] = 8'b10010001;
DRAM[49415] = 8'b10010010;
DRAM[49416] = 8'b10010101;
DRAM[49417] = 8'b10010011;
DRAM[49418] = 8'b10010001;
DRAM[49419] = 8'b10010010;
DRAM[49420] = 8'b10010100;
DRAM[49421] = 8'b10010111;
DRAM[49422] = 8'b10010111;
DRAM[49423] = 8'b10010111;
DRAM[49424] = 8'b10011001;
DRAM[49425] = 8'b10011000;
DRAM[49426] = 8'b10010111;
DRAM[49427] = 8'b10010110;
DRAM[49428] = 8'b10010110;
DRAM[49429] = 8'b10010110;
DRAM[49430] = 8'b10010110;
DRAM[49431] = 8'b10010110;
DRAM[49432] = 8'b10001111;
DRAM[49433] = 8'b10010110;
DRAM[49434] = 8'b10011010;
DRAM[49435] = 8'b10011001;
DRAM[49436] = 8'b10011111;
DRAM[49437] = 8'b10110111;
DRAM[49438] = 8'b11011001;
DRAM[49439] = 8'b11110011;
DRAM[49440] = 8'b11111100;
DRAM[49441] = 8'b11111101;
DRAM[49442] = 8'b11111110;
DRAM[49443] = 8'b11111110;
DRAM[49444] = 8'b11111111;
DRAM[49445] = 8'b11111111;
DRAM[49446] = 8'b11111111;
DRAM[49447] = 8'b11111110;
DRAM[49448] = 8'b11111101;
DRAM[49449] = 8'b11111101;
DRAM[49450] = 8'b11111101;
DRAM[49451] = 8'b11111100;
DRAM[49452] = 8'b11111010;
DRAM[49453] = 8'b11110111;
DRAM[49454] = 8'b11110101;
DRAM[49455] = 8'b11110100;
DRAM[49456] = 8'b11101100;
DRAM[49457] = 8'b11101011;
DRAM[49458] = 8'b11100010;
DRAM[49459] = 8'b11011110;
DRAM[49460] = 8'b11100001;
DRAM[49461] = 8'b11011010;
DRAM[49462] = 8'b11010111;
DRAM[49463] = 8'b11100000;
DRAM[49464] = 8'b11100010;
DRAM[49465] = 8'b11100001;
DRAM[49466] = 8'b11100000;
DRAM[49467] = 8'b11100000;
DRAM[49468] = 8'b11100000;
DRAM[49469] = 8'b11011110;
DRAM[49470] = 8'b11011100;
DRAM[49471] = 8'b11011001;
DRAM[49472] = 8'b11011100;
DRAM[49473] = 8'b11010111;
DRAM[49474] = 8'b11010000;
DRAM[49475] = 8'b11001100;
DRAM[49476] = 8'b11001010;
DRAM[49477] = 8'b11000111;
DRAM[49478] = 8'b11000000;
DRAM[49479] = 8'b10111010;
DRAM[49480] = 8'b10111001;
DRAM[49481] = 8'b10101110;
DRAM[49482] = 8'b10100010;
DRAM[49483] = 8'b10011100;
DRAM[49484] = 8'b10010111;
DRAM[49485] = 8'b10010011;
DRAM[49486] = 8'b10010101;
DRAM[49487] = 8'b10011011;
DRAM[49488] = 8'b10000110;
DRAM[49489] = 8'b10000010;
DRAM[49490] = 8'b10000011;
DRAM[49491] = 8'b10000000;
DRAM[49492] = 8'b1110000;
DRAM[49493] = 8'b1100100;
DRAM[49494] = 8'b1110010;
DRAM[49495] = 8'b10001011;
DRAM[49496] = 8'b10000011;
DRAM[49497] = 8'b1111010;
DRAM[49498] = 8'b1111101;
DRAM[49499] = 8'b10001011;
DRAM[49500] = 8'b10010011;
DRAM[49501] = 8'b10010000;
DRAM[49502] = 8'b10001011;
DRAM[49503] = 8'b10001001;
DRAM[49504] = 8'b10000011;
DRAM[49505] = 8'b10001011;
DRAM[49506] = 8'b1111111;
DRAM[49507] = 8'b1111011;
DRAM[49508] = 8'b1110101;
DRAM[49509] = 8'b1101111;
DRAM[49510] = 8'b1111010;
DRAM[49511] = 8'b1110100;
DRAM[49512] = 8'b1101100;
DRAM[49513] = 8'b1101011;
DRAM[49514] = 8'b1101101;
DRAM[49515] = 8'b1110010;
DRAM[49516] = 8'b1110111;
DRAM[49517] = 8'b1110111;
DRAM[49518] = 8'b1110001;
DRAM[49519] = 8'b1101011;
DRAM[49520] = 8'b1110001;
DRAM[49521] = 8'b1110101;
DRAM[49522] = 8'b1111011;
DRAM[49523] = 8'b1111110;
DRAM[49524] = 8'b10000000;
DRAM[49525] = 8'b10000010;
DRAM[49526] = 8'b10000110;
DRAM[49527] = 8'b10001001;
DRAM[49528] = 8'b1111101;
DRAM[49529] = 8'b1111101;
DRAM[49530] = 8'b10000010;
DRAM[49531] = 8'b10001100;
DRAM[49532] = 8'b10010111;
DRAM[49533] = 8'b10011010;
DRAM[49534] = 8'b10010100;
DRAM[49535] = 8'b10001101;
DRAM[49536] = 8'b10000001;
DRAM[49537] = 8'b10000011;
DRAM[49538] = 8'b10000010;
DRAM[49539] = 8'b1111110;
DRAM[49540] = 8'b1111100;
DRAM[49541] = 8'b1111011;
DRAM[49542] = 8'b1110100;
DRAM[49543] = 8'b1101100;
DRAM[49544] = 8'b1101100;
DRAM[49545] = 8'b1101110;
DRAM[49546] = 8'b1101101;
DRAM[49547] = 8'b1101001;
DRAM[49548] = 8'b1100111;
DRAM[49549] = 8'b1100011;
DRAM[49550] = 8'b1011010;
DRAM[49551] = 8'b1010000;
DRAM[49552] = 8'b1010110;
DRAM[49553] = 8'b1011010;
DRAM[49554] = 8'b1011101;
DRAM[49555] = 8'b1011011;
DRAM[49556] = 8'b1011001;
DRAM[49557] = 8'b1011011;
DRAM[49558] = 8'b1100000;
DRAM[49559] = 8'b1100100;
DRAM[49560] = 8'b1011110;
DRAM[49561] = 8'b1011010;
DRAM[49562] = 8'b1011111;
DRAM[49563] = 8'b1100001;
DRAM[49564] = 8'b1011110;
DRAM[49565] = 8'b1101010;
DRAM[49566] = 8'b1111010;
DRAM[49567] = 8'b1111110;
DRAM[49568] = 8'b1111011;
DRAM[49569] = 8'b10000101;
DRAM[49570] = 8'b10011001;
DRAM[49571] = 8'b10100101;
DRAM[49572] = 8'b10110011;
DRAM[49573] = 8'b10101011;
DRAM[49574] = 8'b10001100;
DRAM[49575] = 8'b10000101;
DRAM[49576] = 8'b10010010;
DRAM[49577] = 8'b10001110;
DRAM[49578] = 8'b10001110;
DRAM[49579] = 8'b10010101;
DRAM[49580] = 8'b10011100;
DRAM[49581] = 8'b10011111;
DRAM[49582] = 8'b10100011;
DRAM[49583] = 8'b10100111;
DRAM[49584] = 8'b10100101;
DRAM[49585] = 8'b10101011;
DRAM[49586] = 8'b10110101;
DRAM[49587] = 8'b11000000;
DRAM[49588] = 8'b11001100;
DRAM[49589] = 8'b11011010;
DRAM[49590] = 8'b11101001;
DRAM[49591] = 8'b11110010;
DRAM[49592] = 8'b11110100;
DRAM[49593] = 8'b11110110;
DRAM[49594] = 8'b11111000;
DRAM[49595] = 8'b11111001;
DRAM[49596] = 8'b11111001;
DRAM[49597] = 8'b11111010;
DRAM[49598] = 8'b11111100;
DRAM[49599] = 8'b11111110;
DRAM[49600] = 8'b11110111;
DRAM[49601] = 8'b11111101;
DRAM[49602] = 8'b11111010;
DRAM[49603] = 8'b11101100;
DRAM[49604] = 8'b11100001;
DRAM[49605] = 8'b11011100;
DRAM[49606] = 8'b11010011;
DRAM[49607] = 8'b11000111;
DRAM[49608] = 8'b10110000;
DRAM[49609] = 8'b10101000;
DRAM[49610] = 8'b10100000;
DRAM[49611] = 8'b10011011;
DRAM[49612] = 8'b10010100;
DRAM[49613] = 8'b10001001;
DRAM[49614] = 8'b10000010;
DRAM[49615] = 8'b10000001;
DRAM[49616] = 8'b1111110;
DRAM[49617] = 8'b1111101;
DRAM[49618] = 8'b1111011;
DRAM[49619] = 8'b1111001;
DRAM[49620] = 8'b1110110;
DRAM[49621] = 8'b1110100;
DRAM[49622] = 8'b1110010;
DRAM[49623] = 8'b1110001;
DRAM[49624] = 8'b1101111;
DRAM[49625] = 8'b1101111;
DRAM[49626] = 8'b1101110;
DRAM[49627] = 8'b1101110;
DRAM[49628] = 8'b1101111;
DRAM[49629] = 8'b1110000;
DRAM[49630] = 8'b1110010;
DRAM[49631] = 8'b1110011;
DRAM[49632] = 8'b1110100;
DRAM[49633] = 8'b1110101;
DRAM[49634] = 8'b1110110;
DRAM[49635] = 8'b1111000;
DRAM[49636] = 8'b1111001;
DRAM[49637] = 8'b1111010;
DRAM[49638] = 8'b1111010;
DRAM[49639] = 8'b1111010;
DRAM[49640] = 8'b1111010;
DRAM[49641] = 8'b1111010;
DRAM[49642] = 8'b1111011;
DRAM[49643] = 8'b1111011;
DRAM[49644] = 8'b1111101;
DRAM[49645] = 8'b1111110;
DRAM[49646] = 8'b10000000;
DRAM[49647] = 8'b10000001;
DRAM[49648] = 8'b10000001;
DRAM[49649] = 8'b10000001;
DRAM[49650] = 8'b10000010;
DRAM[49651] = 8'b10000010;
DRAM[49652] = 8'b10000011;
DRAM[49653] = 8'b10000011;
DRAM[49654] = 8'b10000011;
DRAM[49655] = 8'b10000011;
DRAM[49656] = 8'b10000010;
DRAM[49657] = 8'b10000010;
DRAM[49658] = 8'b10000010;
DRAM[49659] = 8'b10000011;
DRAM[49660] = 8'b10000011;
DRAM[49661] = 8'b10000100;
DRAM[49662] = 8'b10000100;
DRAM[49663] = 8'b10000100;
DRAM[49664] = 8'b10001100;
DRAM[49665] = 8'b10001100;
DRAM[49666] = 8'b10001101;
DRAM[49667] = 8'b10001111;
DRAM[49668] = 8'b10010000;
DRAM[49669] = 8'b10010010;
DRAM[49670] = 8'b10010011;
DRAM[49671] = 8'b10010100;
DRAM[49672] = 8'b10010101;
DRAM[49673] = 8'b10010100;
DRAM[49674] = 8'b10010011;
DRAM[49675] = 8'b10010011;
DRAM[49676] = 8'b10010110;
DRAM[49677] = 8'b10011000;
DRAM[49678] = 8'b10011000;
DRAM[49679] = 8'b10010111;
DRAM[49680] = 8'b10011000;
DRAM[49681] = 8'b10011000;
DRAM[49682] = 8'b10010111;
DRAM[49683] = 8'b10010110;
DRAM[49684] = 8'b10010110;
DRAM[49685] = 8'b10010110;
DRAM[49686] = 8'b10010110;
DRAM[49687] = 8'b10010111;
DRAM[49688] = 8'b10010010;
DRAM[49689] = 8'b10011000;
DRAM[49690] = 8'b10010110;
DRAM[49691] = 8'b10010010;
DRAM[49692] = 8'b10100011;
DRAM[49693] = 8'b11001001;
DRAM[49694] = 8'b11101001;
DRAM[49695] = 8'b11110110;
DRAM[49696] = 8'b11111100;
DRAM[49697] = 8'b11111101;
DRAM[49698] = 8'b11111101;
DRAM[49699] = 8'b11111110;
DRAM[49700] = 8'b11111111;
DRAM[49701] = 8'b11111110;
DRAM[49702] = 8'b11111110;
DRAM[49703] = 8'b11111110;
DRAM[49704] = 8'b11111011;
DRAM[49705] = 8'b11111101;
DRAM[49706] = 8'b11111111;
DRAM[49707] = 8'b11111111;
DRAM[49708] = 8'b11111110;
DRAM[49709] = 8'b11111011;
DRAM[49710] = 8'b11110111;
DRAM[49711] = 8'b11110100;
DRAM[49712] = 8'b11101110;
DRAM[49713] = 8'b11101111;
DRAM[49714] = 8'b11101000;
DRAM[49715] = 8'b11100110;
DRAM[49716] = 8'b11101001;
DRAM[49717] = 8'b11100001;
DRAM[49718] = 8'b11011010;
DRAM[49719] = 8'b11100010;
DRAM[49720] = 8'b11100000;
DRAM[49721] = 8'b11011101;
DRAM[49722] = 8'b11011001;
DRAM[49723] = 8'b11011001;
DRAM[49724] = 8'b11011010;
DRAM[49725] = 8'b11011010;
DRAM[49726] = 8'b11011000;
DRAM[49727] = 8'b11010110;
DRAM[49728] = 8'b11011000;
DRAM[49729] = 8'b11010100;
DRAM[49730] = 8'b11001101;
DRAM[49731] = 8'b11001001;
DRAM[49732] = 8'b11000100;
DRAM[49733] = 8'b10111110;
DRAM[49734] = 8'b10110101;
DRAM[49735] = 8'b10101110;
DRAM[49736] = 8'b10110010;
DRAM[49737] = 8'b10100110;
DRAM[49738] = 8'b10011001;
DRAM[49739] = 8'b10010100;
DRAM[49740] = 8'b10010010;
DRAM[49741] = 8'b10010010;
DRAM[49742] = 8'b10010011;
DRAM[49743] = 8'b10010101;
DRAM[49744] = 8'b10001011;
DRAM[49745] = 8'b10001100;
DRAM[49746] = 8'b10001100;
DRAM[49747] = 8'b10001010;
DRAM[49748] = 8'b10000100;
DRAM[49749] = 8'b10000011;
DRAM[49750] = 8'b10001101;
DRAM[49751] = 8'b10011010;
DRAM[49752] = 8'b10001011;
DRAM[49753] = 8'b1111001;
DRAM[49754] = 8'b1111111;
DRAM[49755] = 8'b10001101;
DRAM[49756] = 8'b10001000;
DRAM[49757] = 8'b10000111;
DRAM[49758] = 8'b10001010;
DRAM[49759] = 8'b10000001;
DRAM[49760] = 8'b1111101;
DRAM[49761] = 8'b10001110;
DRAM[49762] = 8'b10000010;
DRAM[49763] = 8'b1111000;
DRAM[49764] = 8'b1110111;
DRAM[49765] = 8'b1111100;
DRAM[49766] = 8'b1111110;
DRAM[49767] = 8'b1100110;
DRAM[49768] = 8'b1100101;
DRAM[49769] = 8'b1100101;
DRAM[49770] = 8'b1101101;
DRAM[49771] = 8'b1111000;
DRAM[49772] = 8'b1111000;
DRAM[49773] = 8'b1101111;
DRAM[49774] = 8'b1101011;
DRAM[49775] = 8'b1101110;
DRAM[49776] = 8'b1101000;
DRAM[49777] = 8'b1101000;
DRAM[49778] = 8'b1101010;
DRAM[49779] = 8'b1101100;
DRAM[49780] = 8'b1110000;
DRAM[49781] = 8'b1110101;
DRAM[49782] = 8'b1111010;
DRAM[49783] = 8'b1111110;
DRAM[49784] = 8'b1110011;
DRAM[49785] = 8'b1110101;
DRAM[49786] = 8'b1111010;
DRAM[49787] = 8'b10000100;
DRAM[49788] = 8'b10001111;
DRAM[49789] = 8'b10010110;
DRAM[49790] = 8'b10011000;
DRAM[49791] = 8'b10010111;
DRAM[49792] = 8'b10001111;
DRAM[49793] = 8'b10001101;
DRAM[49794] = 8'b10000110;
DRAM[49795] = 8'b10000000;
DRAM[49796] = 8'b1111111;
DRAM[49797] = 8'b10000000;
DRAM[49798] = 8'b1111010;
DRAM[49799] = 8'b1110001;
DRAM[49800] = 8'b1110011;
DRAM[49801] = 8'b1110011;
DRAM[49802] = 8'b1101110;
DRAM[49803] = 8'b1101000;
DRAM[49804] = 8'b1100101;
DRAM[49805] = 8'b1100101;
DRAM[49806] = 8'b1100001;
DRAM[49807] = 8'b1011100;
DRAM[49808] = 8'b1100010;
DRAM[49809] = 8'b1100001;
DRAM[49810] = 8'b1100000;
DRAM[49811] = 8'b1011111;
DRAM[49812] = 8'b1011110;
DRAM[49813] = 8'b1011111;
DRAM[49814] = 8'b1100000;
DRAM[49815] = 8'b1100010;
DRAM[49816] = 8'b1101000;
DRAM[49817] = 8'b1100111;
DRAM[49818] = 8'b1110000;
DRAM[49819] = 8'b1110011;
DRAM[49820] = 8'b1101101;
DRAM[49821] = 8'b1110100;
DRAM[49822] = 8'b10000010;
DRAM[49823] = 8'b10000111;
DRAM[49824] = 8'b10001001;
DRAM[49825] = 8'b10011110;
DRAM[49826] = 8'b10100011;
DRAM[49827] = 8'b10110001;
DRAM[49828] = 8'b10110111;
DRAM[49829] = 8'b10100001;
DRAM[49830] = 8'b10001011;
DRAM[49831] = 8'b1111001;
DRAM[49832] = 8'b10000111;
DRAM[49833] = 8'b10001000;
DRAM[49834] = 8'b10001101;
DRAM[49835] = 8'b10010101;
DRAM[49836] = 8'b10011010;
DRAM[49837] = 8'b10011011;
DRAM[49838] = 8'b10011111;
DRAM[49839] = 8'b10100101;
DRAM[49840] = 8'b10100111;
DRAM[49841] = 8'b10101000;
DRAM[49842] = 8'b10101100;
DRAM[49843] = 8'b10110101;
DRAM[49844] = 8'b11000100;
DRAM[49845] = 8'b11010110;
DRAM[49846] = 8'b11100100;
DRAM[49847] = 8'b11101101;
DRAM[49848] = 8'b11110100;
DRAM[49849] = 8'b11110110;
DRAM[49850] = 8'b11111001;
DRAM[49851] = 8'b11111010;
DRAM[49852] = 8'b11111001;
DRAM[49853] = 8'b11111001;
DRAM[49854] = 8'b11111010;
DRAM[49855] = 8'b11111011;
DRAM[49856] = 8'b11111011;
DRAM[49857] = 8'b11111111;
DRAM[49858] = 8'b11110110;
DRAM[49859] = 8'b11011110;
DRAM[49860] = 8'b11000110;
DRAM[49861] = 8'b10111011;
DRAM[49862] = 8'b10110110;
DRAM[49863] = 8'b10110010;
DRAM[49864] = 8'b10101111;
DRAM[49865] = 8'b10100110;
DRAM[49866] = 8'b10011101;
DRAM[49867] = 8'b10010111;
DRAM[49868] = 8'b10010000;
DRAM[49869] = 8'b10000111;
DRAM[49870] = 8'b10000001;
DRAM[49871] = 8'b10000000;
DRAM[49872] = 8'b1111100;
DRAM[49873] = 8'b1111011;
DRAM[49874] = 8'b1111010;
DRAM[49875] = 8'b1110111;
DRAM[49876] = 8'b1110101;
DRAM[49877] = 8'b1110010;
DRAM[49878] = 8'b1110001;
DRAM[49879] = 8'b1110000;
DRAM[49880] = 8'b1101110;
DRAM[49881] = 8'b1101101;
DRAM[49882] = 8'b1101101;
DRAM[49883] = 8'b1101101;
DRAM[49884] = 8'b1101110;
DRAM[49885] = 8'b1110000;
DRAM[49886] = 8'b1110001;
DRAM[49887] = 8'b1110010;
DRAM[49888] = 8'b1110100;
DRAM[49889] = 8'b1110101;
DRAM[49890] = 8'b1110110;
DRAM[49891] = 8'b1111000;
DRAM[49892] = 8'b1111001;
DRAM[49893] = 8'b1111010;
DRAM[49894] = 8'b1111010;
DRAM[49895] = 8'b1111010;
DRAM[49896] = 8'b1111011;
DRAM[49897] = 8'b1111010;
DRAM[49898] = 8'b1111011;
DRAM[49899] = 8'b1111011;
DRAM[49900] = 8'b1111100;
DRAM[49901] = 8'b1111110;
DRAM[49902] = 8'b1111111;
DRAM[49903] = 8'b10000000;
DRAM[49904] = 8'b1111111;
DRAM[49905] = 8'b1111111;
DRAM[49906] = 8'b10000000;
DRAM[49907] = 8'b10000000;
DRAM[49908] = 8'b10000000;
DRAM[49909] = 8'b10000001;
DRAM[49910] = 8'b10000001;
DRAM[49911] = 8'b10000001;
DRAM[49912] = 8'b1111111;
DRAM[49913] = 8'b10000000;
DRAM[49914] = 8'b10000000;
DRAM[49915] = 8'b10000000;
DRAM[49916] = 8'b10000000;
DRAM[49917] = 8'b10000001;
DRAM[49918] = 8'b10000001;
DRAM[49919] = 8'b10000001;
DRAM[49920] = 8'b10001100;
DRAM[49921] = 8'b10001101;
DRAM[49922] = 8'b10001110;
DRAM[49923] = 8'b10001111;
DRAM[49924] = 8'b10010001;
DRAM[49925] = 8'b10010010;
DRAM[49926] = 8'b10010011;
DRAM[49927] = 8'b10010011;
DRAM[49928] = 8'b10010110;
DRAM[49929] = 8'b10010100;
DRAM[49930] = 8'b10010011;
DRAM[49931] = 8'b10010101;
DRAM[49932] = 8'b10010111;
DRAM[49933] = 8'b10011001;
DRAM[49934] = 8'b10011000;
DRAM[49935] = 8'b10010111;
DRAM[49936] = 8'b10010111;
DRAM[49937] = 8'b10010111;
DRAM[49938] = 8'b10010110;
DRAM[49939] = 8'b10010101;
DRAM[49940] = 8'b10010101;
DRAM[49941] = 8'b10010110;
DRAM[49942] = 8'b10010110;
DRAM[49943] = 8'b10010111;
DRAM[49944] = 8'b10010111;
DRAM[49945] = 8'b10011000;
DRAM[49946] = 8'b10010110;
DRAM[49947] = 8'b10011000;
DRAM[49948] = 8'b10101100;
DRAM[49949] = 8'b11001110;
DRAM[49950] = 8'b11101010;
DRAM[49951] = 8'b11110110;
DRAM[49952] = 8'b11111100;
DRAM[49953] = 8'b11111101;
DRAM[49954] = 8'b11111101;
DRAM[49955] = 8'b11111110;
DRAM[49956] = 8'b11111110;
DRAM[49957] = 8'b11111110;
DRAM[49958] = 8'b11111101;
DRAM[49959] = 8'b11111101;
DRAM[49960] = 8'b11111011;
DRAM[49961] = 8'b11111100;
DRAM[49962] = 8'b11111101;
DRAM[49963] = 8'b11111110;
DRAM[49964] = 8'b11111101;
DRAM[49965] = 8'b11111011;
DRAM[49966] = 8'b11111000;
DRAM[49967] = 8'b11110110;
DRAM[49968] = 8'b11110000;
DRAM[49969] = 8'b11110010;
DRAM[49970] = 8'b11101100;
DRAM[49971] = 8'b11101010;
DRAM[49972] = 8'b11101100;
DRAM[49973] = 8'b11100010;
DRAM[49974] = 8'b11011001;
DRAM[49975] = 8'b11011111;
DRAM[49976] = 8'b11011011;
DRAM[49977] = 8'b11010111;
DRAM[49978] = 8'b11010101;
DRAM[49979] = 8'b11010101;
DRAM[49980] = 8'b11011000;
DRAM[49981] = 8'b11011001;
DRAM[49982] = 8'b11010110;
DRAM[49983] = 8'b11010010;
DRAM[49984] = 8'b11010010;
DRAM[49985] = 8'b11001111;
DRAM[49986] = 8'b11001011;
DRAM[49987] = 8'b11000110;
DRAM[49988] = 8'b11000001;
DRAM[49989] = 8'b10111010;
DRAM[49990] = 8'b10110001;
DRAM[49991] = 8'b10101011;
DRAM[49992] = 8'b10100011;
DRAM[49993] = 8'b10010111;
DRAM[49994] = 8'b10001110;
DRAM[49995] = 8'b10010010;
DRAM[49996] = 8'b10011011;
DRAM[49997] = 8'b10011101;
DRAM[49998] = 8'b10010010;
DRAM[49999] = 8'b10001000;
DRAM[50000] = 8'b10000011;
DRAM[50001] = 8'b10001000;
DRAM[50002] = 8'b10001011;
DRAM[50003] = 8'b10001110;
DRAM[50004] = 8'b10010010;
DRAM[50005] = 8'b10010111;
DRAM[50006] = 8'b10010110;
DRAM[50007] = 8'b10010010;
DRAM[50008] = 8'b10010000;
DRAM[50009] = 8'b1111010;
DRAM[50010] = 8'b10000110;
DRAM[50011] = 8'b10010100;
DRAM[50012] = 8'b10000101;
DRAM[50013] = 8'b10000100;
DRAM[50014] = 8'b10001010;
DRAM[50015] = 8'b1111100;
DRAM[50016] = 8'b1111100;
DRAM[50017] = 8'b10001001;
DRAM[50018] = 8'b1111100;
DRAM[50019] = 8'b1110111;
DRAM[50020] = 8'b1111001;
DRAM[50021] = 8'b1111101;
DRAM[50022] = 8'b1111101;
DRAM[50023] = 8'b1100001;
DRAM[50024] = 8'b1110010;
DRAM[50025] = 8'b1101010;
DRAM[50026] = 8'b1101011;
DRAM[50027] = 8'b1110011;
DRAM[50028] = 8'b1110001;
DRAM[50029] = 8'b1100110;
DRAM[50030] = 8'b1100110;
DRAM[50031] = 8'b1110000;
DRAM[50032] = 8'b1100110;
DRAM[50033] = 8'b1100011;
DRAM[50034] = 8'b1100001;
DRAM[50035] = 8'b1100010;
DRAM[50036] = 8'b1100101;
DRAM[50037] = 8'b1101000;
DRAM[50038] = 8'b1101010;
DRAM[50039] = 8'b1101011;
DRAM[50040] = 8'b1100000;
DRAM[50041] = 8'b1100110;
DRAM[50042] = 8'b1101110;
DRAM[50043] = 8'b1110100;
DRAM[50044] = 8'b1111011;
DRAM[50045] = 8'b10000011;
DRAM[50046] = 8'b10001110;
DRAM[50047] = 8'b10010101;
DRAM[50048] = 8'b10011001;
DRAM[50049] = 8'b10010111;
DRAM[50050] = 8'b10001111;
DRAM[50051] = 8'b10000101;
DRAM[50052] = 8'b10000001;
DRAM[50053] = 8'b10000010;
DRAM[50054] = 8'b10000000;
DRAM[50055] = 8'b1111100;
DRAM[50056] = 8'b1111111;
DRAM[50057] = 8'b1111010;
DRAM[50058] = 8'b1101110;
DRAM[50059] = 8'b1100010;
DRAM[50060] = 8'b1011111;
DRAM[50061] = 8'b1100101;
DRAM[50062] = 8'b1101011;
DRAM[50063] = 8'b1101100;
DRAM[50064] = 8'b1101010;
DRAM[50065] = 8'b1100100;
DRAM[50066] = 8'b1100000;
DRAM[50067] = 8'b1100010;
DRAM[50068] = 8'b1100011;
DRAM[50069] = 8'b1100010;
DRAM[50070] = 8'b1100001;
DRAM[50071] = 8'b1100010;
DRAM[50072] = 8'b1101110;
DRAM[50073] = 8'b1101011;
DRAM[50074] = 8'b1110101;
DRAM[50075] = 8'b1111110;
DRAM[50076] = 8'b1111011;
DRAM[50077] = 8'b10000000;
DRAM[50078] = 8'b10001011;
DRAM[50079] = 8'b10001100;
DRAM[50080] = 8'b10011101;
DRAM[50081] = 8'b10101110;
DRAM[50082] = 8'b10011001;
DRAM[50083] = 8'b10011100;
DRAM[50084] = 8'b10011110;
DRAM[50085] = 8'b10001111;
DRAM[50086] = 8'b10010110;
DRAM[50087] = 8'b10001100;
DRAM[50088] = 8'b10000100;
DRAM[50089] = 8'b10001000;
DRAM[50090] = 8'b10001111;
DRAM[50091] = 8'b10010110;
DRAM[50092] = 8'b10010111;
DRAM[50093] = 8'b10010111;
DRAM[50094] = 8'b10011101;
DRAM[50095] = 8'b10100110;
DRAM[50096] = 8'b10101010;
DRAM[50097] = 8'b10101100;
DRAM[50098] = 8'b10101111;
DRAM[50099] = 8'b10110111;
DRAM[50100] = 8'b11000010;
DRAM[50101] = 8'b11010000;
DRAM[50102] = 8'b11011111;
DRAM[50103] = 8'b11101000;
DRAM[50104] = 8'b11110100;
DRAM[50105] = 8'b11110110;
DRAM[50106] = 8'b11110111;
DRAM[50107] = 8'b11110111;
DRAM[50108] = 8'b11110110;
DRAM[50109] = 8'b11110111;
DRAM[50110] = 8'b11111001;
DRAM[50111] = 8'b11111011;
DRAM[50112] = 8'b11111000;
DRAM[50113] = 8'b11111010;
DRAM[50114] = 8'b11101111;
DRAM[50115] = 8'b11010110;
DRAM[50116] = 8'b10111101;
DRAM[50117] = 8'b10101111;
DRAM[50118] = 8'b10101010;
DRAM[50119] = 8'b10101000;
DRAM[50120] = 8'b10110011;
DRAM[50121] = 8'b10100111;
DRAM[50122] = 8'b10011010;
DRAM[50123] = 8'b10010001;
DRAM[50124] = 8'b10001010;
DRAM[50125] = 8'b10000011;
DRAM[50126] = 8'b10000001;
DRAM[50127] = 8'b10000010;
DRAM[50128] = 8'b1111100;
DRAM[50129] = 8'b1111011;
DRAM[50130] = 8'b1111001;
DRAM[50131] = 8'b1110111;
DRAM[50132] = 8'b1110100;
DRAM[50133] = 8'b1110010;
DRAM[50134] = 8'b1110000;
DRAM[50135] = 8'b1101111;
DRAM[50136] = 8'b1101110;
DRAM[50137] = 8'b1101110;
DRAM[50138] = 8'b1101110;
DRAM[50139] = 8'b1101111;
DRAM[50140] = 8'b1101111;
DRAM[50141] = 8'b1110000;
DRAM[50142] = 8'b1110001;
DRAM[50143] = 8'b1110010;
DRAM[50144] = 8'b1110011;
DRAM[50145] = 8'b1110100;
DRAM[50146] = 8'b1110110;
DRAM[50147] = 8'b1110111;
DRAM[50148] = 8'b1111001;
DRAM[50149] = 8'b1111001;
DRAM[50150] = 8'b1111010;
DRAM[50151] = 8'b1111010;
DRAM[50152] = 8'b1111011;
DRAM[50153] = 8'b1111011;
DRAM[50154] = 8'b1111011;
DRAM[50155] = 8'b1111011;
DRAM[50156] = 8'b1111100;
DRAM[50157] = 8'b1111101;
DRAM[50158] = 8'b1111111;
DRAM[50159] = 8'b1111111;
DRAM[50160] = 8'b1111111;
DRAM[50161] = 8'b1111111;
DRAM[50162] = 8'b1111111;
DRAM[50163] = 8'b1111111;
DRAM[50164] = 8'b1111111;
DRAM[50165] = 8'b1111111;
DRAM[50166] = 8'b1111111;
DRAM[50167] = 8'b1111111;
DRAM[50168] = 8'b1111110;
DRAM[50169] = 8'b1111110;
DRAM[50170] = 8'b1111110;
DRAM[50171] = 8'b1111111;
DRAM[50172] = 8'b1111111;
DRAM[50173] = 8'b1111111;
DRAM[50174] = 8'b1111111;
DRAM[50175] = 8'b1111111;
DRAM[50176] = 8'b10001100;
DRAM[50177] = 8'b10001100;
DRAM[50178] = 8'b10001101;
DRAM[50179] = 8'b10001110;
DRAM[50180] = 8'b10001111;
DRAM[50181] = 8'b10010000;
DRAM[50182] = 8'b10010001;
DRAM[50183] = 8'b10010001;
DRAM[50184] = 8'b10010101;
DRAM[50185] = 8'b10010100;
DRAM[50186] = 8'b10010100;
DRAM[50187] = 8'b10010101;
DRAM[50188] = 8'b10011000;
DRAM[50189] = 8'b10011001;
DRAM[50190] = 8'b10011000;
DRAM[50191] = 8'b10010111;
DRAM[50192] = 8'b10010110;
DRAM[50193] = 8'b10010110;
DRAM[50194] = 8'b10010101;
DRAM[50195] = 8'b10010101;
DRAM[50196] = 8'b10010101;
DRAM[50197] = 8'b10010110;
DRAM[50198] = 8'b10010110;
DRAM[50199] = 8'b10010111;
DRAM[50200] = 8'b10011000;
DRAM[50201] = 8'b10010100;
DRAM[50202] = 8'b10011000;
DRAM[50203] = 8'b10101000;
DRAM[50204] = 8'b10111011;
DRAM[50205] = 8'b11001110;
DRAM[50206] = 8'b11100101;
DRAM[50207] = 8'b11111001;
DRAM[50208] = 8'b11111100;
DRAM[50209] = 8'b11111101;
DRAM[50210] = 8'b11111101;
DRAM[50211] = 8'b11111110;
DRAM[50212] = 8'b11111110;
DRAM[50213] = 8'b11111101;
DRAM[50214] = 8'b11111100;
DRAM[50215] = 8'b11111100;
DRAM[50216] = 8'b11111100;
DRAM[50217] = 8'b11111100;
DRAM[50218] = 8'b11111010;
DRAM[50219] = 8'b11111001;
DRAM[50220] = 8'b11111000;
DRAM[50221] = 8'b11111000;
DRAM[50222] = 8'b11110111;
DRAM[50223] = 8'b11110111;
DRAM[50224] = 8'b11101110;
DRAM[50225] = 8'b11101111;
DRAM[50226] = 8'b11101001;
DRAM[50227] = 8'b11100110;
DRAM[50228] = 8'b11100110;
DRAM[50229] = 8'b11011011;
DRAM[50230] = 8'b11010001;
DRAM[50231] = 8'b11010111;
DRAM[50232] = 8'b11011011;
DRAM[50233] = 8'b11011010;
DRAM[50234] = 8'b11011011;
DRAM[50235] = 8'b11011101;
DRAM[50236] = 8'b11100000;
DRAM[50237] = 8'b11011111;
DRAM[50238] = 8'b11011010;
DRAM[50239] = 8'b11010110;
DRAM[50240] = 8'b11010010;
DRAM[50241] = 8'b11001111;
DRAM[50242] = 8'b11001011;
DRAM[50243] = 8'b11000110;
DRAM[50244] = 8'b11000000;
DRAM[50245] = 8'b10111000;
DRAM[50246] = 8'b10110000;
DRAM[50247] = 8'b10101011;
DRAM[50248] = 8'b10011001;
DRAM[50249] = 8'b10010110;
DRAM[50250] = 8'b10010101;
DRAM[50251] = 8'b10010111;
DRAM[50252] = 8'b10011100;
DRAM[50253] = 8'b10011100;
DRAM[50254] = 8'b10010100;
DRAM[50255] = 8'b10001011;
DRAM[50256] = 8'b10000100;
DRAM[50257] = 8'b10010010;
DRAM[50258] = 8'b10011011;
DRAM[50259] = 8'b10010111;
DRAM[50260] = 8'b10010001;
DRAM[50261] = 8'b10010010;
DRAM[50262] = 8'b10010101;
DRAM[50263] = 8'b10010101;
DRAM[50264] = 8'b10001111;
DRAM[50265] = 8'b1111011;
DRAM[50266] = 8'b10001011;
DRAM[50267] = 8'b10011010;
DRAM[50268] = 8'b10000111;
DRAM[50269] = 8'b10000010;
DRAM[50270] = 8'b10001000;
DRAM[50271] = 8'b1111001;
DRAM[50272] = 8'b10000011;
DRAM[50273] = 8'b10000011;
DRAM[50274] = 8'b1110110;
DRAM[50275] = 8'b1111100;
DRAM[50276] = 8'b1111111;
DRAM[50277] = 8'b1111000;
DRAM[50278] = 8'b1111000;
DRAM[50279] = 8'b1101010;
DRAM[50280] = 8'b1110110;
DRAM[50281] = 8'b1101010;
DRAM[50282] = 8'b1100110;
DRAM[50283] = 8'b1101101;
DRAM[50284] = 8'b1101100;
DRAM[50285] = 8'b1100001;
DRAM[50286] = 8'b1100000;
DRAM[50287] = 8'b1101001;
DRAM[50288] = 8'b1100111;
DRAM[50289] = 8'b1100110;
DRAM[50290] = 8'b1100101;
DRAM[50291] = 8'b1100101;
DRAM[50292] = 8'b1100101;
DRAM[50293] = 8'b1100101;
DRAM[50294] = 8'b1100011;
DRAM[50295] = 8'b1100001;
DRAM[50296] = 8'b1010101;
DRAM[50297] = 8'b1011110;
DRAM[50298] = 8'b1100110;
DRAM[50299] = 8'b1100110;
DRAM[50300] = 8'b1100100;
DRAM[50301] = 8'b1101001;
DRAM[50302] = 8'b1110110;
DRAM[50303] = 8'b10000011;
DRAM[50304] = 8'b10001100;
DRAM[50305] = 8'b10010100;
DRAM[50306] = 8'b10011000;
DRAM[50307] = 8'b10010010;
DRAM[50308] = 8'b10001100;
DRAM[50309] = 8'b10001010;
DRAM[50310] = 8'b10001010;
DRAM[50311] = 8'b10001000;
DRAM[50312] = 8'b10000101;
DRAM[50313] = 8'b10000001;
DRAM[50314] = 8'b1110110;
DRAM[50315] = 8'b1101010;
DRAM[50316] = 8'b1100111;
DRAM[50317] = 8'b1101101;
DRAM[50318] = 8'b1110100;
DRAM[50319] = 8'b1110111;
DRAM[50320] = 8'b1110001;
DRAM[50321] = 8'b1101001;
DRAM[50322] = 8'b1100101;
DRAM[50323] = 8'b1101001;
DRAM[50324] = 8'b1101100;
DRAM[50325] = 8'b1101011;
DRAM[50326] = 8'b1101010;
DRAM[50327] = 8'b1101011;
DRAM[50328] = 8'b1110011;
DRAM[50329] = 8'b1101100;
DRAM[50330] = 8'b1110110;
DRAM[50331] = 8'b10000111;
DRAM[50332] = 8'b10001100;
DRAM[50333] = 8'b10010011;
DRAM[50334] = 8'b10011001;
DRAM[50335] = 8'b10010111;
DRAM[50336] = 8'b10011001;
DRAM[50337] = 8'b10100111;
DRAM[50338] = 8'b10001000;
DRAM[50339] = 8'b10000000;
DRAM[50340] = 8'b10000000;
DRAM[50341] = 8'b1111011;
DRAM[50342] = 8'b10010001;
DRAM[50343] = 8'b10010010;
DRAM[50344] = 8'b10000100;
DRAM[50345] = 8'b10001000;
DRAM[50346] = 8'b10001110;
DRAM[50347] = 8'b10010100;
DRAM[50348] = 8'b10010100;
DRAM[50349] = 8'b10010100;
DRAM[50350] = 8'b10011100;
DRAM[50351] = 8'b10100110;
DRAM[50352] = 8'b10100101;
DRAM[50353] = 8'b10101100;
DRAM[50354] = 8'b10110101;
DRAM[50355] = 8'b10111011;
DRAM[50356] = 8'b11000001;
DRAM[50357] = 8'b11001011;
DRAM[50358] = 8'b11011010;
DRAM[50359] = 8'b11100110;
DRAM[50360] = 8'b11110100;
DRAM[50361] = 8'b11110100;
DRAM[50362] = 8'b11110100;
DRAM[50363] = 8'b11110010;
DRAM[50364] = 8'b11110010;
DRAM[50365] = 8'b11110100;
DRAM[50366] = 8'b11111000;
DRAM[50367] = 8'b11111100;
DRAM[50368] = 8'b11110100;
DRAM[50369] = 8'b11110011;
DRAM[50370] = 8'b11101010;
DRAM[50371] = 8'b11011010;
DRAM[50372] = 8'b11001010;
DRAM[50373] = 8'b10111110;
DRAM[50374] = 8'b10110110;
DRAM[50375] = 8'b10110000;
DRAM[50376] = 8'b10101000;
DRAM[50377] = 8'b10011111;
DRAM[50378] = 8'b10010110;
DRAM[50379] = 8'b10010001;
DRAM[50380] = 8'b10001011;
DRAM[50381] = 8'b10000011;
DRAM[50382] = 8'b1111111;
DRAM[50383] = 8'b1111111;
DRAM[50384] = 8'b1111101;
DRAM[50385] = 8'b1111100;
DRAM[50386] = 8'b1111010;
DRAM[50387] = 8'b1111000;
DRAM[50388] = 8'b1110101;
DRAM[50389] = 8'b1110011;
DRAM[50390] = 8'b1110001;
DRAM[50391] = 8'b1110000;
DRAM[50392] = 8'b1101110;
DRAM[50393] = 8'b1101111;
DRAM[50394] = 8'b1110000;
DRAM[50395] = 8'b1110001;
DRAM[50396] = 8'b1110001;
DRAM[50397] = 8'b1110010;
DRAM[50398] = 8'b1110010;
DRAM[50399] = 8'b1110010;
DRAM[50400] = 8'b1110011;
DRAM[50401] = 8'b1110100;
DRAM[50402] = 8'b1110101;
DRAM[50403] = 8'b1110111;
DRAM[50404] = 8'b1111000;
DRAM[50405] = 8'b1111001;
DRAM[50406] = 8'b1111001;
DRAM[50407] = 8'b1111001;
DRAM[50408] = 8'b1111011;
DRAM[50409] = 8'b1111011;
DRAM[50410] = 8'b1111010;
DRAM[50411] = 8'b1111011;
DRAM[50412] = 8'b1111011;
DRAM[50413] = 8'b1111100;
DRAM[50414] = 8'b1111110;
DRAM[50415] = 8'b1111110;
DRAM[50416] = 8'b1111111;
DRAM[50417] = 8'b1111111;
DRAM[50418] = 8'b1111111;
DRAM[50419] = 8'b1111111;
DRAM[50420] = 8'b1111111;
DRAM[50421] = 8'b1111111;
DRAM[50422] = 8'b1111111;
DRAM[50423] = 8'b1111111;
DRAM[50424] = 8'b1111110;
DRAM[50425] = 8'b1111110;
DRAM[50426] = 8'b1111110;
DRAM[50427] = 8'b1111101;
DRAM[50428] = 8'b1111101;
DRAM[50429] = 8'b1111101;
DRAM[50430] = 8'b1111101;
DRAM[50431] = 8'b1111101;
DRAM[50432] = 8'b10001011;
DRAM[50433] = 8'b10001011;
DRAM[50434] = 8'b10001100;
DRAM[50435] = 8'b10001101;
DRAM[50436] = 8'b10001110;
DRAM[50437] = 8'b10001111;
DRAM[50438] = 8'b10001111;
DRAM[50439] = 8'b10010000;
DRAM[50440] = 8'b10010100;
DRAM[50441] = 8'b10010011;
DRAM[50442] = 8'b10010011;
DRAM[50443] = 8'b10010101;
DRAM[50444] = 8'b10011000;
DRAM[50445] = 8'b10011000;
DRAM[50446] = 8'b10010111;
DRAM[50447] = 8'b10010101;
DRAM[50448] = 8'b10010101;
DRAM[50449] = 8'b10010101;
DRAM[50450] = 8'b10010101;
DRAM[50451] = 8'b10010100;
DRAM[50452] = 8'b10010101;
DRAM[50453] = 8'b10010110;
DRAM[50454] = 8'b10010110;
DRAM[50455] = 8'b10010111;
DRAM[50456] = 8'b10010101;
DRAM[50457] = 8'b10010010;
DRAM[50458] = 8'b10011110;
DRAM[50459] = 8'b10110110;
DRAM[50460] = 8'b11001010;
DRAM[50461] = 8'b11010110;
DRAM[50462] = 8'b11101010;
DRAM[50463] = 8'b11111111;
DRAM[50464] = 8'b11111100;
DRAM[50465] = 8'b11111101;
DRAM[50466] = 8'b11111101;
DRAM[50467] = 8'b11111101;
DRAM[50468] = 8'b11111101;
DRAM[50469] = 8'b11111100;
DRAM[50470] = 8'b11111011;
DRAM[50471] = 8'b11111011;
DRAM[50472] = 8'b11111101;
DRAM[50473] = 8'b11111011;
DRAM[50474] = 8'b11111001;
DRAM[50475] = 8'b11110111;
DRAM[50476] = 8'b11110101;
DRAM[50477] = 8'b11110101;
DRAM[50478] = 8'b11110101;
DRAM[50479] = 8'b11110110;
DRAM[50480] = 8'b11110000;
DRAM[50481] = 8'b11110000;
DRAM[50482] = 8'b11100111;
DRAM[50483] = 8'b11100011;
DRAM[50484] = 8'b11100011;
DRAM[50485] = 8'b11011001;
DRAM[50486] = 8'b11010001;
DRAM[50487] = 8'b11010111;
DRAM[50488] = 8'b11011001;
DRAM[50489] = 8'b11011011;
DRAM[50490] = 8'b11011110;
DRAM[50491] = 8'b11100000;
DRAM[50492] = 8'b11011111;
DRAM[50493] = 8'b11011011;
DRAM[50494] = 8'b11010111;
DRAM[50495] = 8'b11010101;
DRAM[50496] = 8'b11001101;
DRAM[50497] = 8'b11001011;
DRAM[50498] = 8'b11000110;
DRAM[50499] = 8'b10111111;
DRAM[50500] = 8'b10110111;
DRAM[50501] = 8'b10101111;
DRAM[50502] = 8'b10101000;
DRAM[50503] = 8'b10100100;
DRAM[50504] = 8'b10011101;
DRAM[50505] = 8'b10100101;
DRAM[50506] = 8'b10101000;
DRAM[50507] = 8'b10100000;
DRAM[50508] = 8'b10010110;
DRAM[50509] = 8'b10010100;
DRAM[50510] = 8'b10011010;
DRAM[50511] = 8'b10011110;
DRAM[50512] = 8'b10101011;
DRAM[50513] = 8'b10100111;
DRAM[50514] = 8'b10100000;
DRAM[50515] = 8'b10011011;
DRAM[50516] = 8'b10011100;
DRAM[50517] = 8'b10011110;
DRAM[50518] = 8'b10011011;
DRAM[50519] = 8'b10010101;
DRAM[50520] = 8'b10001101;
DRAM[50521] = 8'b10000010;
DRAM[50522] = 8'b10001110;
DRAM[50523] = 8'b10011001;
DRAM[50524] = 8'b10001011;
DRAM[50525] = 8'b10000001;
DRAM[50526] = 8'b10000001;
DRAM[50527] = 8'b1111010;
DRAM[50528] = 8'b10001010;
DRAM[50529] = 8'b10000100;
DRAM[50530] = 8'b1111000;
DRAM[50531] = 8'b10000101;
DRAM[50532] = 8'b10000100;
DRAM[50533] = 8'b1110001;
DRAM[50534] = 8'b1110011;
DRAM[50535] = 8'b1110001;
DRAM[50536] = 8'b1101000;
DRAM[50537] = 8'b1100011;
DRAM[50538] = 8'b1100101;
DRAM[50539] = 8'b1101100;
DRAM[50540] = 8'b1101011;
DRAM[50541] = 8'b1100010;
DRAM[50542] = 8'b1011101;
DRAM[50543] = 8'b1011111;
DRAM[50544] = 8'b1100011;
DRAM[50545] = 8'b1100100;
DRAM[50546] = 8'b1100101;
DRAM[50547] = 8'b1100101;
DRAM[50548] = 8'b1100100;
DRAM[50549] = 8'b1100001;
DRAM[50550] = 8'b1011110;
DRAM[50551] = 8'b1011100;
DRAM[50552] = 8'b1011001;
DRAM[50553] = 8'b1011111;
DRAM[50554] = 8'b1100011;
DRAM[50555] = 8'b1011111;
DRAM[50556] = 8'b1011000;
DRAM[50557] = 8'b1011000;
DRAM[50558] = 8'b1100010;
DRAM[50559] = 8'b1101100;
DRAM[50560] = 8'b1110001;
DRAM[50561] = 8'b10000011;
DRAM[50562] = 8'b10010100;
DRAM[50563] = 8'b10011000;
DRAM[50564] = 8'b10010100;
DRAM[50565] = 8'b10010001;
DRAM[50566] = 8'b10001111;
DRAM[50567] = 8'b10001101;
DRAM[50568] = 8'b10000100;
DRAM[50569] = 8'b10000111;
DRAM[50570] = 8'b10000110;
DRAM[50571] = 8'b10000000;
DRAM[50572] = 8'b1111100;
DRAM[50573] = 8'b1111101;
DRAM[50574] = 8'b1111100;
DRAM[50575] = 8'b1111010;
DRAM[50576] = 8'b1110100;
DRAM[50577] = 8'b1101100;
DRAM[50578] = 8'b1101001;
DRAM[50579] = 8'b1101111;
DRAM[50580] = 8'b1110011;
DRAM[50581] = 8'b1110000;
DRAM[50582] = 8'b1110000;
DRAM[50583] = 8'b1110100;
DRAM[50584] = 8'b1111110;
DRAM[50585] = 8'b1110011;
DRAM[50586] = 8'b1111100;
DRAM[50587] = 8'b10010001;
DRAM[50588] = 8'b10011001;
DRAM[50589] = 8'b10011110;
DRAM[50590] = 8'b10100010;
DRAM[50591] = 8'b10011110;
DRAM[50592] = 8'b10000110;
DRAM[50593] = 8'b10010110;
DRAM[50594] = 8'b10001010;
DRAM[50595] = 8'b1111110;
DRAM[50596] = 8'b1111100;
DRAM[50597] = 8'b1111010;
DRAM[50598] = 8'b10000100;
DRAM[50599] = 8'b10001000;
DRAM[50600] = 8'b10001111;
DRAM[50601] = 8'b10010000;
DRAM[50602] = 8'b10010011;
DRAM[50603] = 8'b10010100;
DRAM[50604] = 8'b10010001;
DRAM[50605] = 8'b10001101;
DRAM[50606] = 8'b10010001;
DRAM[50607] = 8'b10011000;
DRAM[50608] = 8'b10011011;
DRAM[50609] = 8'b10100101;
DRAM[50610] = 8'b10110010;
DRAM[50611] = 8'b10111010;
DRAM[50612] = 8'b10111111;
DRAM[50613] = 8'b11001000;
DRAM[50614] = 8'b11010111;
DRAM[50615] = 8'b11100011;
DRAM[50616] = 8'b11101111;
DRAM[50617] = 8'b11110000;
DRAM[50618] = 8'b11110001;
DRAM[50619] = 8'b11110000;
DRAM[50620] = 8'b11110000;
DRAM[50621] = 8'b11110011;
DRAM[50622] = 8'b11110111;
DRAM[50623] = 8'b11111010;
DRAM[50624] = 8'b11110111;
DRAM[50625] = 8'b11110100;
DRAM[50626] = 8'b11101100;
DRAM[50627] = 8'b11100001;
DRAM[50628] = 8'b11010011;
DRAM[50629] = 8'b11000011;
DRAM[50630] = 8'b10110100;
DRAM[50631] = 8'b10101010;
DRAM[50632] = 8'b10011000;
DRAM[50633] = 8'b10010100;
DRAM[50634] = 8'b10010011;
DRAM[50635] = 8'b10010100;
DRAM[50636] = 8'b10010000;
DRAM[50637] = 8'b10000110;
DRAM[50638] = 8'b1111100;
DRAM[50639] = 8'b1111001;
DRAM[50640] = 8'b1111100;
DRAM[50641] = 8'b1111011;
DRAM[50642] = 8'b1111010;
DRAM[50643] = 8'b1110111;
DRAM[50644] = 8'b1110101;
DRAM[50645] = 8'b1110010;
DRAM[50646] = 8'b1110001;
DRAM[50647] = 8'b1110000;
DRAM[50648] = 8'b1101110;
DRAM[50649] = 8'b1101111;
DRAM[50650] = 8'b1110000;
DRAM[50651] = 8'b1110010;
DRAM[50652] = 8'b1110011;
DRAM[50653] = 8'b1110011;
DRAM[50654] = 8'b1110011;
DRAM[50655] = 8'b1110010;
DRAM[50656] = 8'b1110010;
DRAM[50657] = 8'b1110011;
DRAM[50658] = 8'b1110101;
DRAM[50659] = 8'b1110111;
DRAM[50660] = 8'b1111000;
DRAM[50661] = 8'b1111001;
DRAM[50662] = 8'b1111001;
DRAM[50663] = 8'b1111001;
DRAM[50664] = 8'b1111011;
DRAM[50665] = 8'b1111011;
DRAM[50666] = 8'b1111010;
DRAM[50667] = 8'b1111010;
DRAM[50668] = 8'b1111011;
DRAM[50669] = 8'b1111100;
DRAM[50670] = 8'b1111101;
DRAM[50671] = 8'b1111101;
DRAM[50672] = 8'b1111111;
DRAM[50673] = 8'b1111111;
DRAM[50674] = 8'b1111110;
DRAM[50675] = 8'b1111110;
DRAM[50676] = 8'b1111110;
DRAM[50677] = 8'b1111101;
DRAM[50678] = 8'b1111101;
DRAM[50679] = 8'b1111101;
DRAM[50680] = 8'b1111101;
DRAM[50681] = 8'b1111100;
DRAM[50682] = 8'b1111100;
DRAM[50683] = 8'b1111100;
DRAM[50684] = 8'b1111100;
DRAM[50685] = 8'b1111011;
DRAM[50686] = 8'b1111011;
DRAM[50687] = 8'b1111011;
DRAM[50688] = 8'b10001011;
DRAM[50689] = 8'b10001100;
DRAM[50690] = 8'b10001100;
DRAM[50691] = 8'b10001101;
DRAM[50692] = 8'b10001110;
DRAM[50693] = 8'b10001110;
DRAM[50694] = 8'b10001111;
DRAM[50695] = 8'b10001111;
DRAM[50696] = 8'b10010010;
DRAM[50697] = 8'b10010010;
DRAM[50698] = 8'b10010011;
DRAM[50699] = 8'b10010101;
DRAM[50700] = 8'b10010111;
DRAM[50701] = 8'b10011000;
DRAM[50702] = 8'b10010110;
DRAM[50703] = 8'b10010100;
DRAM[50704] = 8'b10010101;
DRAM[50705] = 8'b10010100;
DRAM[50706] = 8'b10010100;
DRAM[50707] = 8'b10010100;
DRAM[50708] = 8'b10010101;
DRAM[50709] = 8'b10010101;
DRAM[50710] = 8'b10010110;
DRAM[50711] = 8'b10010111;
DRAM[50712] = 8'b10010111;
DRAM[50713] = 8'b10011011;
DRAM[50714] = 8'b10101000;
DRAM[50715] = 8'b10111101;
DRAM[50716] = 8'b11010100;
DRAM[50717] = 8'b11100111;
DRAM[50718] = 8'b11110110;
DRAM[50719] = 8'b11111111;
DRAM[50720] = 8'b11111101;
DRAM[50721] = 8'b11111101;
DRAM[50722] = 8'b11111101;
DRAM[50723] = 8'b11111101;
DRAM[50724] = 8'b11111101;
DRAM[50725] = 8'b11111100;
DRAM[50726] = 8'b11111011;
DRAM[50727] = 8'b11111010;
DRAM[50728] = 8'b11111100;
DRAM[50729] = 8'b11111011;
DRAM[50730] = 8'b11111010;
DRAM[50731] = 8'b11111001;
DRAM[50732] = 8'b11110111;
DRAM[50733] = 8'b11110101;
DRAM[50734] = 8'b11110011;
DRAM[50735] = 8'b11110010;
DRAM[50736] = 8'b11110001;
DRAM[50737] = 8'b11110000;
DRAM[50738] = 8'b11100110;
DRAM[50739] = 8'b11100001;
DRAM[50740] = 8'b11100010;
DRAM[50741] = 8'b11011010;
DRAM[50742] = 8'b11010110;
DRAM[50743] = 8'b11011110;
DRAM[50744] = 8'b11010111;
DRAM[50745] = 8'b11011011;
DRAM[50746] = 8'b11011101;
DRAM[50747] = 8'b11011010;
DRAM[50748] = 8'b11010011;
DRAM[50749] = 8'b11001110;
DRAM[50750] = 8'b11001101;
DRAM[50751] = 8'b11001110;
DRAM[50752] = 8'b11000110;
DRAM[50753] = 8'b11000100;
DRAM[50754] = 8'b11000000;
DRAM[50755] = 8'b10111001;
DRAM[50756] = 8'b10110010;
DRAM[50757] = 8'b10101011;
DRAM[50758] = 8'b10100111;
DRAM[50759] = 8'b10100101;
DRAM[50760] = 8'b10101100;
DRAM[50761] = 8'b10110001;
DRAM[50762] = 8'b10110000;
DRAM[50763] = 8'b10100110;
DRAM[50764] = 8'b10011110;
DRAM[50765] = 8'b10100001;
DRAM[50766] = 8'b10100111;
DRAM[50767] = 8'b10101010;
DRAM[50768] = 8'b10110101;
DRAM[50769] = 8'b10100010;
DRAM[50770] = 8'b10010001;
DRAM[50771] = 8'b10010011;
DRAM[50772] = 8'b10011110;
DRAM[50773] = 8'b10100000;
DRAM[50774] = 8'b10010100;
DRAM[50775] = 8'b10000111;
DRAM[50776] = 8'b10010010;
DRAM[50777] = 8'b10001111;
DRAM[50778] = 8'b10010011;
DRAM[50779] = 8'b10011000;
DRAM[50780] = 8'b10001111;
DRAM[50781] = 8'b10000001;
DRAM[50782] = 8'b1111101;
DRAM[50783] = 8'b10000000;
DRAM[50784] = 8'b10001010;
DRAM[50785] = 8'b10001010;
DRAM[50786] = 8'b10000001;
DRAM[50787] = 8'b10001011;
DRAM[50788] = 8'b10000010;
DRAM[50789] = 8'b1101011;
DRAM[50790] = 8'b1101110;
DRAM[50791] = 8'b1101110;
DRAM[50792] = 8'b1011111;
DRAM[50793] = 8'b1100101;
DRAM[50794] = 8'b1101100;
DRAM[50795] = 8'b1101110;
DRAM[50796] = 8'b1101001;
DRAM[50797] = 8'b1100010;
DRAM[50798] = 8'b1011111;
DRAM[50799] = 8'b1011110;
DRAM[50800] = 8'b1100001;
DRAM[50801] = 8'b1100100;
DRAM[50802] = 8'b1100110;
DRAM[50803] = 8'b1100100;
DRAM[50804] = 8'b1011111;
DRAM[50805] = 8'b1011011;
DRAM[50806] = 8'b1011010;
DRAM[50807] = 8'b1011010;
DRAM[50808] = 8'b1011110;
DRAM[50809] = 8'b1011110;
DRAM[50810] = 8'b1011100;
DRAM[50811] = 8'b1011010;
DRAM[50812] = 8'b1011001;
DRAM[50813] = 8'b1011001;
DRAM[50814] = 8'b1011010;
DRAM[50815] = 8'b1011100;
DRAM[50816] = 8'b1100010;
DRAM[50817] = 8'b1110001;
DRAM[50818] = 8'b1111111;
DRAM[50819] = 8'b10000101;
DRAM[50820] = 8'b10000110;
DRAM[50821] = 8'b10001001;
DRAM[50822] = 8'b10001010;
DRAM[50823] = 8'b10001010;
DRAM[50824] = 8'b10000100;
DRAM[50825] = 8'b10001011;
DRAM[50826] = 8'b10010000;
DRAM[50827] = 8'b10001101;
DRAM[50828] = 8'b10001001;
DRAM[50829] = 8'b10000111;
DRAM[50830] = 8'b10000011;
DRAM[50831] = 8'b1111110;
DRAM[50832] = 8'b1111011;
DRAM[50833] = 8'b1110011;
DRAM[50834] = 8'b1110001;
DRAM[50835] = 8'b1111001;
DRAM[50836] = 8'b1111011;
DRAM[50837] = 8'b1110110;
DRAM[50838] = 8'b1111000;
DRAM[50839] = 8'b1111111;
DRAM[50840] = 8'b10001101;
DRAM[50841] = 8'b10000001;
DRAM[50842] = 8'b10001000;
DRAM[50843] = 8'b10010111;
DRAM[50844] = 8'b10010111;
DRAM[50845] = 8'b10010100;
DRAM[50846] = 8'b10010100;
DRAM[50847] = 8'b10010010;
DRAM[50848] = 8'b1111010;
DRAM[50849] = 8'b10001011;
DRAM[50850] = 8'b10010110;
DRAM[50851] = 8'b10000110;
DRAM[50852] = 8'b10000011;
DRAM[50853] = 8'b10000110;
DRAM[50854] = 8'b1111111;
DRAM[50855] = 8'b10001000;
DRAM[50856] = 8'b10010011;
DRAM[50857] = 8'b10010011;
DRAM[50858] = 8'b10010110;
DRAM[50859] = 8'b10011001;
DRAM[50860] = 8'b10010110;
DRAM[50861] = 8'b10010000;
DRAM[50862] = 8'b10001111;
DRAM[50863] = 8'b10010011;
DRAM[50864] = 8'b10011100;
DRAM[50865] = 8'b10100011;
DRAM[50866] = 8'b10101100;
DRAM[50867] = 8'b10110100;
DRAM[50868] = 8'b10111100;
DRAM[50869] = 8'b11000110;
DRAM[50870] = 8'b11010011;
DRAM[50871] = 8'b11011100;
DRAM[50872] = 8'b11100111;
DRAM[50873] = 8'b11101011;
DRAM[50874] = 8'b11101111;
DRAM[50875] = 8'b11110001;
DRAM[50876] = 8'b11110010;
DRAM[50877] = 8'b11110011;
DRAM[50878] = 8'b11110100;
DRAM[50879] = 8'b11110110;
DRAM[50880] = 8'b11111000;
DRAM[50881] = 8'b11110101;
DRAM[50882] = 8'b11101111;
DRAM[50883] = 8'b11100101;
DRAM[50884] = 8'b11010101;
DRAM[50885] = 8'b11000001;
DRAM[50886] = 8'b10101111;
DRAM[50887] = 8'b10100101;
DRAM[50888] = 8'b10011101;
DRAM[50889] = 8'b10011000;
DRAM[50890] = 8'b10010101;
DRAM[50891] = 8'b10010100;
DRAM[50892] = 8'b10001111;
DRAM[50893] = 8'b10000101;
DRAM[50894] = 8'b1111100;
DRAM[50895] = 8'b1111001;
DRAM[50896] = 8'b1111011;
DRAM[50897] = 8'b1111010;
DRAM[50898] = 8'b1111000;
DRAM[50899] = 8'b1110110;
DRAM[50900] = 8'b1110011;
DRAM[50901] = 8'b1110001;
DRAM[50902] = 8'b1101111;
DRAM[50903] = 8'b1101110;
DRAM[50904] = 8'b1101101;
DRAM[50905] = 8'b1101110;
DRAM[50906] = 8'b1110000;
DRAM[50907] = 8'b1110001;
DRAM[50908] = 8'b1110010;
DRAM[50909] = 8'b1110010;
DRAM[50910] = 8'b1110001;
DRAM[50911] = 8'b1110001;
DRAM[50912] = 8'b1110010;
DRAM[50913] = 8'b1110011;
DRAM[50914] = 8'b1110101;
DRAM[50915] = 8'b1110110;
DRAM[50916] = 8'b1111000;
DRAM[50917] = 8'b1111000;
DRAM[50918] = 8'b1111000;
DRAM[50919] = 8'b1111000;
DRAM[50920] = 8'b1111011;
DRAM[50921] = 8'b1111011;
DRAM[50922] = 8'b1111010;
DRAM[50923] = 8'b1111010;
DRAM[50924] = 8'b1111010;
DRAM[50925] = 8'b1111011;
DRAM[50926] = 8'b1111100;
DRAM[50927] = 8'b1111101;
DRAM[50928] = 8'b1111101;
DRAM[50929] = 8'b1111101;
DRAM[50930] = 8'b1111100;
DRAM[50931] = 8'b1111100;
DRAM[50932] = 8'b1111011;
DRAM[50933] = 8'b1111011;
DRAM[50934] = 8'b1111011;
DRAM[50935] = 8'b1111011;
DRAM[50936] = 8'b1111010;
DRAM[50937] = 8'b1111010;
DRAM[50938] = 8'b1111010;
DRAM[50939] = 8'b1111001;
DRAM[50940] = 8'b1111001;
DRAM[50941] = 8'b1111000;
DRAM[50942] = 8'b1111000;
DRAM[50943] = 8'b1111000;
DRAM[50944] = 8'b10001100;
DRAM[50945] = 8'b10001100;
DRAM[50946] = 8'b10001101;
DRAM[50947] = 8'b10001110;
DRAM[50948] = 8'b10001110;
DRAM[50949] = 8'b10001111;
DRAM[50950] = 8'b10001111;
DRAM[50951] = 8'b10010000;
DRAM[50952] = 8'b10010001;
DRAM[50953] = 8'b10010001;
DRAM[50954] = 8'b10010010;
DRAM[50955] = 8'b10010100;
DRAM[50956] = 8'b10010111;
DRAM[50957] = 8'b10010111;
DRAM[50958] = 8'b10010101;
DRAM[50959] = 8'b10010011;
DRAM[50960] = 8'b10010100;
DRAM[50961] = 8'b10010100;
DRAM[50962] = 8'b10010100;
DRAM[50963] = 8'b10010100;
DRAM[50964] = 8'b10010100;
DRAM[50965] = 8'b10010101;
DRAM[50966] = 8'b10010111;
DRAM[50967] = 8'b10010111;
DRAM[50968] = 8'b10011101;
DRAM[50969] = 8'b10100111;
DRAM[50970] = 8'b10110001;
DRAM[50971] = 8'b10111110;
DRAM[50972] = 8'b11010111;
DRAM[50973] = 8'b11110100;
DRAM[50974] = 8'b11111111;
DRAM[50975] = 8'b11111010;
DRAM[50976] = 8'b11111101;
DRAM[50977] = 8'b11111101;
DRAM[50978] = 8'b11111101;
DRAM[50979] = 8'b11111101;
DRAM[50980] = 8'b11111101;
DRAM[50981] = 8'b11111011;
DRAM[50982] = 8'b11111010;
DRAM[50983] = 8'b11111010;
DRAM[50984] = 8'b11111011;
DRAM[50985] = 8'b11111100;
DRAM[50986] = 8'b11111100;
DRAM[50987] = 8'b11111100;
DRAM[50988] = 8'b11111010;
DRAM[50989] = 8'b11110110;
DRAM[50990] = 8'b11110010;
DRAM[50991] = 8'b11101111;
DRAM[50992] = 8'b11101101;
DRAM[50993] = 8'b11101011;
DRAM[50994] = 8'b11100000;
DRAM[50995] = 8'b11011011;
DRAM[50996] = 8'b11011101;
DRAM[50997] = 8'b11011000;
DRAM[50998] = 8'b11010110;
DRAM[50999] = 8'b11100000;
DRAM[51000] = 8'b11011010;
DRAM[51001] = 8'b11011101;
DRAM[51002] = 8'b11011101;
DRAM[51003] = 8'b11010110;
DRAM[51004] = 8'b11001100;
DRAM[51005] = 8'b11000110;
DRAM[51006] = 8'b11000111;
DRAM[51007] = 8'b11001010;
DRAM[51008] = 8'b11000100;
DRAM[51009] = 8'b11000011;
DRAM[51010] = 8'b11000001;
DRAM[51011] = 8'b10111100;
DRAM[51012] = 8'b10110110;
DRAM[51013] = 8'b10110011;
DRAM[51014] = 8'b10110001;
DRAM[51015] = 8'b10110001;
DRAM[51016] = 8'b10111000;
DRAM[51017] = 8'b10110011;
DRAM[51018] = 8'b10101011;
DRAM[51019] = 8'b10101000;
DRAM[51020] = 8'b10110001;
DRAM[51021] = 8'b10111010;
DRAM[51022] = 8'b10110100;
DRAM[51023] = 8'b10101000;
DRAM[51024] = 8'b10100100;
DRAM[51025] = 8'b10100000;
DRAM[51026] = 8'b10100000;
DRAM[51027] = 8'b10100100;
DRAM[51028] = 8'b10100001;
DRAM[51029] = 8'b10010111;
DRAM[51030] = 8'b10010010;
DRAM[51031] = 8'b10010100;
DRAM[51032] = 8'b10011001;
DRAM[51033] = 8'b10011011;
DRAM[51034] = 8'b10011000;
DRAM[51035] = 8'b10010111;
DRAM[51036] = 8'b10010011;
DRAM[51037] = 8'b10000011;
DRAM[51038] = 8'b1111100;
DRAM[51039] = 8'b10000111;
DRAM[51040] = 8'b10000101;
DRAM[51041] = 8'b10001110;
DRAM[51042] = 8'b10001001;
DRAM[51043] = 8'b10001100;
DRAM[51044] = 8'b1111101;
DRAM[51045] = 8'b1100110;
DRAM[51046] = 8'b1101000;
DRAM[51047] = 8'b1100101;
DRAM[51048] = 8'b1100010;
DRAM[51049] = 8'b1101110;
DRAM[51050] = 8'b1110110;
DRAM[51051] = 8'b1101111;
DRAM[51052] = 8'b1100100;
DRAM[51053] = 8'b1100000;
DRAM[51054] = 8'b1100011;
DRAM[51055] = 8'b1100101;
DRAM[51056] = 8'b1101001;
DRAM[51057] = 8'b1101100;
DRAM[51058] = 8'b1101101;
DRAM[51059] = 8'b1101000;
DRAM[51060] = 8'b1100000;
DRAM[51061] = 8'b1011010;
DRAM[51062] = 8'b1011011;
DRAM[51063] = 8'b1011101;
DRAM[51064] = 8'b1011111;
DRAM[51065] = 8'b1011000;
DRAM[51066] = 8'b1010011;
DRAM[51067] = 8'b1010110;
DRAM[51068] = 8'b1011101;
DRAM[51069] = 8'b1100000;
DRAM[51070] = 8'b1011100;
DRAM[51071] = 8'b1010110;
DRAM[51072] = 8'b1100011;
DRAM[51073] = 8'b1100111;
DRAM[51074] = 8'b1101001;
DRAM[51075] = 8'b1101010;
DRAM[51076] = 8'b1101111;
DRAM[51077] = 8'b1111010;
DRAM[51078] = 8'b10000010;
DRAM[51079] = 8'b10000100;
DRAM[51080] = 8'b10001000;
DRAM[51081] = 8'b10001110;
DRAM[51082] = 8'b10010001;
DRAM[51083] = 8'b10001110;
DRAM[51084] = 8'b10001001;
DRAM[51085] = 8'b10001000;
DRAM[51086] = 8'b10000110;
DRAM[51087] = 8'b10000100;
DRAM[51088] = 8'b10000110;
DRAM[51089] = 8'b1111111;
DRAM[51090] = 8'b1111110;
DRAM[51091] = 8'b10000101;
DRAM[51092] = 8'b10000110;
DRAM[51093] = 8'b10000000;
DRAM[51094] = 8'b10000010;
DRAM[51095] = 8'b10001011;
DRAM[51096] = 8'b10011000;
DRAM[51097] = 8'b10001100;
DRAM[51098] = 8'b10010001;
DRAM[51099] = 8'b10011000;
DRAM[51100] = 8'b10001101;
DRAM[51101] = 8'b10000001;
DRAM[51102] = 8'b1111111;
DRAM[51103] = 8'b1111101;
DRAM[51104] = 8'b1110111;
DRAM[51105] = 8'b10000101;
DRAM[51106] = 8'b10011010;
DRAM[51107] = 8'b10000100;
DRAM[51108] = 8'b10000010;
DRAM[51109] = 8'b10001110;
DRAM[51110] = 8'b10000000;
DRAM[51111] = 8'b10010001;
DRAM[51112] = 8'b10000101;
DRAM[51113] = 8'b10001000;
DRAM[51114] = 8'b10010010;
DRAM[51115] = 8'b10011100;
DRAM[51116] = 8'b10100000;
DRAM[51117] = 8'b10011111;
DRAM[51118] = 8'b10011111;
DRAM[51119] = 8'b10100010;
DRAM[51120] = 8'b10100100;
DRAM[51121] = 8'b10100101;
DRAM[51122] = 8'b10101001;
DRAM[51123] = 8'b10110000;
DRAM[51124] = 8'b10111010;
DRAM[51125] = 8'b11000110;
DRAM[51126] = 8'b11010000;
DRAM[51127] = 8'b11010101;
DRAM[51128] = 8'b11100001;
DRAM[51129] = 8'b11100111;
DRAM[51130] = 8'b11101110;
DRAM[51131] = 8'b11110011;
DRAM[51132] = 8'b11110101;
DRAM[51133] = 8'b11110100;
DRAM[51134] = 8'b11110010;
DRAM[51135] = 8'b11110010;
DRAM[51136] = 8'b11110000;
DRAM[51137] = 8'b11110000;
DRAM[51138] = 8'b11101111;
DRAM[51139] = 8'b11101001;
DRAM[51140] = 8'b11011010;
DRAM[51141] = 8'b11001000;
DRAM[51142] = 8'b10111010;
DRAM[51143] = 8'b10110100;
DRAM[51144] = 8'b10110000;
DRAM[51145] = 8'b10100101;
DRAM[51146] = 8'b10011001;
DRAM[51147] = 8'b10010001;
DRAM[51148] = 8'b10001010;
DRAM[51149] = 8'b10000010;
DRAM[51150] = 8'b1111111;
DRAM[51151] = 8'b10000000;
DRAM[51152] = 8'b1111001;
DRAM[51153] = 8'b1111000;
DRAM[51154] = 8'b1110110;
DRAM[51155] = 8'b1110100;
DRAM[51156] = 8'b1110010;
DRAM[51157] = 8'b1101111;
DRAM[51158] = 8'b1101110;
DRAM[51159] = 8'b1101101;
DRAM[51160] = 8'b1101011;
DRAM[51161] = 8'b1101101;
DRAM[51162] = 8'b1101110;
DRAM[51163] = 8'b1110000;
DRAM[51164] = 8'b1110001;
DRAM[51165] = 8'b1110001;
DRAM[51166] = 8'b1110000;
DRAM[51167] = 8'b1101111;
DRAM[51168] = 8'b1110010;
DRAM[51169] = 8'b1110011;
DRAM[51170] = 8'b1110101;
DRAM[51171] = 8'b1110110;
DRAM[51172] = 8'b1110111;
DRAM[51173] = 8'b1111000;
DRAM[51174] = 8'b1111000;
DRAM[51175] = 8'b1111000;
DRAM[51176] = 8'b1111011;
DRAM[51177] = 8'b1111011;
DRAM[51178] = 8'b1111010;
DRAM[51179] = 8'b1111010;
DRAM[51180] = 8'b1111010;
DRAM[51181] = 8'b1111011;
DRAM[51182] = 8'b1111100;
DRAM[51183] = 8'b1111100;
DRAM[51184] = 8'b1111011;
DRAM[51185] = 8'b1111011;
DRAM[51186] = 8'b1111011;
DRAM[51187] = 8'b1111010;
DRAM[51188] = 8'b1111010;
DRAM[51189] = 8'b1111001;
DRAM[51190] = 8'b1111001;
DRAM[51191] = 8'b1111000;
DRAM[51192] = 8'b1111000;
DRAM[51193] = 8'b1111000;
DRAM[51194] = 8'b1111000;
DRAM[51195] = 8'b1110111;
DRAM[51196] = 8'b1110110;
DRAM[51197] = 8'b1110110;
DRAM[51198] = 8'b1110110;
DRAM[51199] = 8'b1110101;
DRAM[51200] = 8'b10001011;
DRAM[51201] = 8'b10001011;
DRAM[51202] = 8'b10001011;
DRAM[51203] = 8'b10001011;
DRAM[51204] = 8'b10001101;
DRAM[51205] = 8'b10010000;
DRAM[51206] = 8'b10010010;
DRAM[51207] = 8'b10010100;
DRAM[51208] = 8'b10010100;
DRAM[51209] = 8'b10010100;
DRAM[51210] = 8'b10010100;
DRAM[51211] = 8'b10010101;
DRAM[51212] = 8'b10010101;
DRAM[51213] = 8'b10010110;
DRAM[51214] = 8'b10010110;
DRAM[51215] = 8'b10010110;
DRAM[51216] = 8'b10010100;
DRAM[51217] = 8'b10010100;
DRAM[51218] = 8'b10010100;
DRAM[51219] = 8'b10010011;
DRAM[51220] = 8'b10010011;
DRAM[51221] = 8'b10010101;
DRAM[51222] = 8'b10011010;
DRAM[51223] = 8'b10011110;
DRAM[51224] = 8'b10100111;
DRAM[51225] = 8'b10101001;
DRAM[51226] = 8'b10110101;
DRAM[51227] = 8'b11001110;
DRAM[51228] = 8'b11101010;
DRAM[51229] = 8'b11111010;
DRAM[51230] = 8'b11111110;
DRAM[51231] = 8'b11111101;
DRAM[51232] = 8'b11111011;
DRAM[51233] = 8'b11111100;
DRAM[51234] = 8'b11111110;
DRAM[51235] = 8'b11111111;
DRAM[51236] = 8'b11111111;
DRAM[51237] = 8'b11111110;
DRAM[51238] = 8'b11111100;
DRAM[51239] = 8'b11111011;
DRAM[51240] = 8'b11111100;
DRAM[51241] = 8'b11111011;
DRAM[51242] = 8'b11111001;
DRAM[51243] = 8'b11110111;
DRAM[51244] = 8'b11110110;
DRAM[51245] = 8'b11110011;
DRAM[51246] = 8'b11101110;
DRAM[51247] = 8'b11101011;
DRAM[51248] = 8'b11101010;
DRAM[51249] = 8'b11100110;
DRAM[51250] = 8'b11100001;
DRAM[51251] = 8'b11011100;
DRAM[51252] = 8'b11011001;
DRAM[51253] = 8'b11010110;
DRAM[51254] = 8'b11010010;
DRAM[51255] = 8'b11001111;
DRAM[51256] = 8'b11000100;
DRAM[51257] = 8'b11000111;
DRAM[51258] = 8'b11000101;
DRAM[51259] = 8'b11000000;
DRAM[51260] = 8'b11000001;
DRAM[51261] = 8'b11000101;
DRAM[51262] = 8'b11000011;
DRAM[51263] = 8'b10111100;
DRAM[51264] = 8'b10111110;
DRAM[51265] = 8'b10111111;
DRAM[51266] = 8'b11000001;
DRAM[51267] = 8'b11000011;
DRAM[51268] = 8'b11000001;
DRAM[51269] = 8'b11000000;
DRAM[51270] = 8'b11001000;
DRAM[51271] = 8'b11010011;
DRAM[51272] = 8'b10100011;
DRAM[51273] = 8'b10101011;
DRAM[51274] = 8'b10110000;
DRAM[51275] = 8'b10110001;
DRAM[51276] = 8'b10110111;
DRAM[51277] = 8'b10111110;
DRAM[51278] = 8'b10111001;
DRAM[51279] = 8'b10101101;
DRAM[51280] = 8'b10101010;
DRAM[51281] = 8'b10100111;
DRAM[51282] = 8'b10100100;
DRAM[51283] = 8'b10100000;
DRAM[51284] = 8'b10011011;
DRAM[51285] = 8'b10010101;
DRAM[51286] = 8'b10001110;
DRAM[51287] = 8'b10001001;
DRAM[51288] = 8'b10010000;
DRAM[51289] = 8'b10010110;
DRAM[51290] = 8'b10011011;
DRAM[51291] = 8'b10011011;
DRAM[51292] = 8'b10010001;
DRAM[51293] = 8'b10001010;
DRAM[51294] = 8'b10001010;
DRAM[51295] = 8'b10001111;
DRAM[51296] = 8'b10001110;
DRAM[51297] = 8'b10001000;
DRAM[51298] = 8'b10001011;
DRAM[51299] = 8'b10000101;
DRAM[51300] = 8'b1101101;
DRAM[51301] = 8'b1100000;
DRAM[51302] = 8'b1100101;
DRAM[51303] = 8'b1101010;
DRAM[51304] = 8'b1100111;
DRAM[51305] = 8'b1101110;
DRAM[51306] = 8'b1110000;
DRAM[51307] = 8'b1101010;
DRAM[51308] = 8'b1101001;
DRAM[51309] = 8'b1101101;
DRAM[51310] = 8'b1101010;
DRAM[51311] = 8'b1100010;
DRAM[51312] = 8'b1101010;
DRAM[51313] = 8'b1100011;
DRAM[51314] = 8'b1011100;
DRAM[51315] = 8'b1011111;
DRAM[51316] = 8'b1100000;
DRAM[51317] = 8'b1010010;
DRAM[51318] = 8'b1010001;
DRAM[51319] = 8'b1100101;
DRAM[51320] = 8'b1100000;
DRAM[51321] = 8'b1011110;
DRAM[51322] = 8'b1011100;
DRAM[51323] = 8'b1011101;
DRAM[51324] = 8'b1011110;
DRAM[51325] = 8'b1011101;
DRAM[51326] = 8'b1011001;
DRAM[51327] = 8'b1010100;
DRAM[51328] = 8'b1010110;
DRAM[51329] = 8'b1100110;
DRAM[51330] = 8'b1011101;
DRAM[51331] = 8'b1011001;
DRAM[51332] = 8'b1011100;
DRAM[51333] = 8'b1100100;
DRAM[51334] = 8'b1110000;
DRAM[51335] = 8'b1100010;
DRAM[51336] = 8'b1111101;
DRAM[51337] = 8'b1111100;
DRAM[51338] = 8'b1111111;
DRAM[51339] = 8'b10000011;
DRAM[51340] = 8'b10000011;
DRAM[51341] = 8'b10000010;
DRAM[51342] = 8'b10000110;
DRAM[51343] = 8'b10001011;
DRAM[51344] = 8'b10000100;
DRAM[51345] = 8'b10000100;
DRAM[51346] = 8'b10000100;
DRAM[51347] = 8'b10000110;
DRAM[51348] = 8'b10001011;
DRAM[51349] = 8'b10001011;
DRAM[51350] = 8'b10000101;
DRAM[51351] = 8'b1111101;
DRAM[51352] = 8'b10010001;
DRAM[51353] = 8'b10000011;
DRAM[51354] = 8'b1110111;
DRAM[51355] = 8'b1110100;
DRAM[51356] = 8'b1110011;
DRAM[51357] = 8'b1110000;
DRAM[51358] = 8'b1110010;
DRAM[51359] = 8'b1111000;
DRAM[51360] = 8'b10000010;
DRAM[51361] = 8'b1111110;
DRAM[51362] = 8'b10000111;
DRAM[51363] = 8'b10011010;
DRAM[51364] = 8'b10011011;
DRAM[51365] = 8'b10001101;
DRAM[51366] = 8'b10000111;
DRAM[51367] = 8'b10001111;
DRAM[51368] = 8'b10010000;
DRAM[51369] = 8'b10001011;
DRAM[51370] = 8'b10001001;
DRAM[51371] = 8'b10010010;
DRAM[51372] = 8'b10011111;
DRAM[51373] = 8'b10100110;
DRAM[51374] = 8'b10100001;
DRAM[51375] = 8'b10011010;
DRAM[51376] = 8'b10100011;
DRAM[51377] = 8'b10100100;
DRAM[51378] = 8'b10101010;
DRAM[51379] = 8'b10110101;
DRAM[51380] = 8'b10111111;
DRAM[51381] = 8'b11001000;
DRAM[51382] = 8'b11010100;
DRAM[51383] = 8'b11011111;
DRAM[51384] = 8'b11011101;
DRAM[51385] = 8'b11100100;
DRAM[51386] = 8'b11101010;
DRAM[51387] = 8'b11101011;
DRAM[51388] = 8'b11101001;
DRAM[51389] = 8'b11101010;
DRAM[51390] = 8'b11110000;
DRAM[51391] = 8'b11110110;
DRAM[51392] = 8'b11110100;
DRAM[51393] = 8'b11110100;
DRAM[51394] = 8'b11110010;
DRAM[51395] = 8'b11101001;
DRAM[51396] = 8'b11011011;
DRAM[51397] = 8'b11001011;
DRAM[51398] = 8'b10111111;
DRAM[51399] = 8'b10111000;
DRAM[51400] = 8'b10100111;
DRAM[51401] = 8'b10011010;
DRAM[51402] = 8'b10001100;
DRAM[51403] = 8'b10000101;
DRAM[51404] = 8'b10000010;
DRAM[51405] = 8'b1111110;
DRAM[51406] = 8'b1111110;
DRAM[51407] = 8'b10000000;
DRAM[51408] = 8'b1111100;
DRAM[51409] = 8'b1111010;
DRAM[51410] = 8'b1110111;
DRAM[51411] = 8'b1110101;
DRAM[51412] = 8'b1110110;
DRAM[51413] = 8'b1110101;
DRAM[51414] = 8'b1110100;
DRAM[51415] = 8'b1110010;
DRAM[51416] = 8'b1101111;
DRAM[51417] = 8'b1101111;
DRAM[51418] = 8'b1101111;
DRAM[51419] = 8'b1110001;
DRAM[51420] = 8'b1110011;
DRAM[51421] = 8'b1110100;
DRAM[51422] = 8'b1110011;
DRAM[51423] = 8'b1110001;
DRAM[51424] = 8'b1110010;
DRAM[51425] = 8'b1110010;
DRAM[51426] = 8'b1110011;
DRAM[51427] = 8'b1110100;
DRAM[51428] = 8'b1110110;
DRAM[51429] = 8'b1110111;
DRAM[51430] = 8'b1111000;
DRAM[51431] = 8'b1111000;
DRAM[51432] = 8'b1111001;
DRAM[51433] = 8'b1111001;
DRAM[51434] = 8'b1111001;
DRAM[51435] = 8'b1111001;
DRAM[51436] = 8'b1111001;
DRAM[51437] = 8'b1111001;
DRAM[51438] = 8'b1111001;
DRAM[51439] = 8'b1111001;
DRAM[51440] = 8'b1111001;
DRAM[51441] = 8'b1111001;
DRAM[51442] = 8'b1111000;
DRAM[51443] = 8'b1111000;
DRAM[51444] = 8'b1110111;
DRAM[51445] = 8'b1110110;
DRAM[51446] = 8'b1110101;
DRAM[51447] = 8'b1110101;
DRAM[51448] = 8'b1110110;
DRAM[51449] = 8'b1110101;
DRAM[51450] = 8'b1110100;
DRAM[51451] = 8'b1110011;
DRAM[51452] = 8'b1110100;
DRAM[51453] = 8'b1110101;
DRAM[51454] = 8'b1110111;
DRAM[51455] = 8'b1111000;
DRAM[51456] = 8'b10001011;
DRAM[51457] = 8'b10001011;
DRAM[51458] = 8'b10001011;
DRAM[51459] = 8'b10001100;
DRAM[51460] = 8'b10001110;
DRAM[51461] = 8'b10010000;
DRAM[51462] = 8'b10010010;
DRAM[51463] = 8'b10010100;
DRAM[51464] = 8'b10010100;
DRAM[51465] = 8'b10010100;
DRAM[51466] = 8'b10010100;
DRAM[51467] = 8'b10010101;
DRAM[51468] = 8'b10010101;
DRAM[51469] = 8'b10010110;
DRAM[51470] = 8'b10010110;
DRAM[51471] = 8'b10010110;
DRAM[51472] = 8'b10010011;
DRAM[51473] = 8'b10010100;
DRAM[51474] = 8'b10010100;
DRAM[51475] = 8'b10010100;
DRAM[51476] = 8'b10010101;
DRAM[51477] = 8'b10011000;
DRAM[51478] = 8'b10011110;
DRAM[51479] = 8'b10100010;
DRAM[51480] = 8'b10101100;
DRAM[51481] = 8'b10110001;
DRAM[51482] = 8'b10111111;
DRAM[51483] = 8'b11010111;
DRAM[51484] = 8'b11101110;
DRAM[51485] = 8'b11111100;
DRAM[51486] = 8'b11111101;
DRAM[51487] = 8'b11111011;
DRAM[51488] = 8'b11111100;
DRAM[51489] = 8'b11111101;
DRAM[51490] = 8'b11111110;
DRAM[51491] = 8'b11111110;
DRAM[51492] = 8'b11111101;
DRAM[51493] = 8'b11111011;
DRAM[51494] = 8'b11111010;
DRAM[51495] = 8'b11111001;
DRAM[51496] = 8'b11111010;
DRAM[51497] = 8'b11111000;
DRAM[51498] = 8'b11110110;
DRAM[51499] = 8'b11110101;
DRAM[51500] = 8'b11110011;
DRAM[51501] = 8'b11110000;
DRAM[51502] = 8'b11101011;
DRAM[51503] = 8'b11100111;
DRAM[51504] = 8'b11011101;
DRAM[51505] = 8'b11011011;
DRAM[51506] = 8'b11011010;
DRAM[51507] = 8'b11011010;
DRAM[51508] = 8'b11011011;
DRAM[51509] = 8'b11011100;
DRAM[51510] = 8'b11011011;
DRAM[51511] = 8'b11011001;
DRAM[51512] = 8'b11000111;
DRAM[51513] = 8'b11001010;
DRAM[51514] = 8'b11001010;
DRAM[51515] = 8'b11000100;
DRAM[51516] = 8'b11000010;
DRAM[51517] = 8'b11000101;
DRAM[51518] = 8'b11000100;
DRAM[51519] = 8'b11000001;
DRAM[51520] = 8'b10111100;
DRAM[51521] = 8'b10111100;
DRAM[51522] = 8'b11000000;
DRAM[51523] = 8'b11000111;
DRAM[51524] = 8'b11000101;
DRAM[51525] = 8'b10111100;
DRAM[51526] = 8'b10110010;
DRAM[51527] = 8'b10101110;
DRAM[51528] = 8'b10101101;
DRAM[51529] = 8'b10111000;
DRAM[51530] = 8'b10111110;
DRAM[51531] = 8'b10111000;
DRAM[51532] = 8'b10101110;
DRAM[51533] = 8'b10101010;
DRAM[51534] = 8'b10101101;
DRAM[51535] = 8'b10110000;
DRAM[51536] = 8'b10101101;
DRAM[51537] = 8'b10101011;
DRAM[51538] = 8'b10101000;
DRAM[51539] = 8'b10100100;
DRAM[51540] = 8'b10100000;
DRAM[51541] = 8'b10011010;
DRAM[51542] = 8'b10010011;
DRAM[51543] = 8'b10001101;
DRAM[51544] = 8'b10001101;
DRAM[51545] = 8'b10010111;
DRAM[51546] = 8'b10010001;
DRAM[51547] = 8'b10100001;
DRAM[51548] = 8'b10001111;
DRAM[51549] = 8'b10010111;
DRAM[51550] = 8'b10001010;
DRAM[51551] = 8'b10001111;
DRAM[51552] = 8'b10000100;
DRAM[51553] = 8'b10000001;
DRAM[51554] = 8'b10000110;
DRAM[51555] = 8'b1111101;
DRAM[51556] = 8'b1100011;
DRAM[51557] = 8'b1011010;
DRAM[51558] = 8'b1100111;
DRAM[51559] = 8'b1110011;
DRAM[51560] = 8'b1100111;
DRAM[51561] = 8'b1101010;
DRAM[51562] = 8'b1101011;
DRAM[51563] = 8'b1101010;
DRAM[51564] = 8'b1101100;
DRAM[51565] = 8'b1101110;
DRAM[51566] = 8'b1101011;
DRAM[51567] = 8'b1100101;
DRAM[51568] = 8'b1100111;
DRAM[51569] = 8'b1100101;
DRAM[51570] = 8'b1011110;
DRAM[51571] = 8'b1011110;
DRAM[51572] = 8'b1011111;
DRAM[51573] = 8'b1010110;
DRAM[51574] = 8'b1010101;
DRAM[51575] = 8'b1100101;
DRAM[51576] = 8'b1011110;
DRAM[51577] = 8'b1011101;
DRAM[51578] = 8'b1011100;
DRAM[51579] = 8'b1011110;
DRAM[51580] = 8'b1100001;
DRAM[51581] = 8'b1011111;
DRAM[51582] = 8'b1011010;
DRAM[51583] = 8'b1010101;
DRAM[51584] = 8'b1011011;
DRAM[51585] = 8'b1101001;
DRAM[51586] = 8'b1011110;
DRAM[51587] = 8'b1010111;
DRAM[51588] = 8'b1010110;
DRAM[51589] = 8'b1011011;
DRAM[51590] = 8'b1100101;
DRAM[51591] = 8'b1010110;
DRAM[51592] = 8'b1101100;
DRAM[51593] = 8'b1101000;
DRAM[51594] = 8'b1101000;
DRAM[51595] = 8'b1101100;
DRAM[51596] = 8'b1101111;
DRAM[51597] = 8'b1110000;
DRAM[51598] = 8'b1110100;
DRAM[51599] = 8'b1111001;
DRAM[51600] = 8'b1111001;
DRAM[51601] = 8'b10000010;
DRAM[51602] = 8'b10000001;
DRAM[51603] = 8'b1111001;
DRAM[51604] = 8'b1111010;
DRAM[51605] = 8'b10000100;
DRAM[51606] = 8'b10000011;
DRAM[51607] = 8'b1111001;
DRAM[51608] = 8'b1111100;
DRAM[51609] = 8'b1110110;
DRAM[51610] = 8'b1110001;
DRAM[51611] = 8'b1110001;
DRAM[51612] = 8'b1110010;
DRAM[51613] = 8'b1110100;
DRAM[51614] = 8'b1110111;
DRAM[51615] = 8'b1111010;
DRAM[51616] = 8'b10000000;
DRAM[51617] = 8'b1111011;
DRAM[51618] = 8'b10000001;
DRAM[51619] = 8'b10001111;
DRAM[51620] = 8'b10010101;
DRAM[51621] = 8'b10001110;
DRAM[51622] = 8'b10001000;
DRAM[51623] = 8'b10001000;
DRAM[51624] = 8'b10010010;
DRAM[51625] = 8'b10001111;
DRAM[51626] = 8'b10001101;
DRAM[51627] = 8'b10010011;
DRAM[51628] = 8'b10011101;
DRAM[51629] = 8'b10100010;
DRAM[51630] = 8'b10100001;
DRAM[51631] = 8'b10011101;
DRAM[51632] = 8'b10100000;
DRAM[51633] = 8'b10100001;
DRAM[51634] = 8'b10101000;
DRAM[51635] = 8'b10110010;
DRAM[51636] = 8'b10111011;
DRAM[51637] = 8'b11000010;
DRAM[51638] = 8'b11001100;
DRAM[51639] = 8'b11010110;
DRAM[51640] = 8'b11100101;
DRAM[51641] = 8'b11101000;
DRAM[51642] = 8'b11101001;
DRAM[51643] = 8'b11100110;
DRAM[51644] = 8'b11100011;
DRAM[51645] = 8'b11100100;
DRAM[51646] = 8'b11101011;
DRAM[51647] = 8'b11110010;
DRAM[51648] = 8'b11111001;
DRAM[51649] = 8'b11110101;
DRAM[51650] = 8'b11101100;
DRAM[51651] = 8'b11011110;
DRAM[51652] = 8'b11001110;
DRAM[51653] = 8'b10111101;
DRAM[51654] = 8'b10110001;
DRAM[51655] = 8'b10101010;
DRAM[51656] = 8'b10100100;
DRAM[51657] = 8'b10011001;
DRAM[51658] = 8'b10001110;
DRAM[51659] = 8'b10001010;
DRAM[51660] = 8'b10000110;
DRAM[51661] = 8'b10000001;
DRAM[51662] = 8'b1111110;
DRAM[51663] = 8'b1111110;
DRAM[51664] = 8'b1111101;
DRAM[51665] = 8'b1111010;
DRAM[51666] = 8'b1110111;
DRAM[51667] = 8'b1110100;
DRAM[51668] = 8'b1110100;
DRAM[51669] = 8'b1110011;
DRAM[51670] = 8'b1110001;
DRAM[51671] = 8'b1101111;
DRAM[51672] = 8'b1101111;
DRAM[51673] = 8'b1101110;
DRAM[51674] = 8'b1101110;
DRAM[51675] = 8'b1110000;
DRAM[51676] = 8'b1110010;
DRAM[51677] = 8'b1110011;
DRAM[51678] = 8'b1110010;
DRAM[51679] = 8'b1110001;
DRAM[51680] = 8'b1110001;
DRAM[51681] = 8'b1110010;
DRAM[51682] = 8'b1110011;
DRAM[51683] = 8'b1110100;
DRAM[51684] = 8'b1110110;
DRAM[51685] = 8'b1110111;
DRAM[51686] = 8'b1111000;
DRAM[51687] = 8'b1111001;
DRAM[51688] = 8'b1111001;
DRAM[51689] = 8'b1111001;
DRAM[51690] = 8'b1111001;
DRAM[51691] = 8'b1111001;
DRAM[51692] = 8'b1111001;
DRAM[51693] = 8'b1111001;
DRAM[51694] = 8'b1111001;
DRAM[51695] = 8'b1111001;
DRAM[51696] = 8'b1110111;
DRAM[51697] = 8'b1110111;
DRAM[51698] = 8'b1110111;
DRAM[51699] = 8'b1110110;
DRAM[51700] = 8'b1110101;
DRAM[51701] = 8'b1110100;
DRAM[51702] = 8'b1110100;
DRAM[51703] = 8'b1110011;
DRAM[51704] = 8'b1110101;
DRAM[51705] = 8'b1110100;
DRAM[51706] = 8'b1110100;
DRAM[51707] = 8'b1110011;
DRAM[51708] = 8'b1110100;
DRAM[51709] = 8'b1110101;
DRAM[51710] = 8'b1110110;
DRAM[51711] = 8'b1110111;
DRAM[51712] = 8'b10001100;
DRAM[51713] = 8'b10001100;
DRAM[51714] = 8'b10001100;
DRAM[51715] = 8'b10001101;
DRAM[51716] = 8'b10001111;
DRAM[51717] = 8'b10010001;
DRAM[51718] = 8'b10010011;
DRAM[51719] = 8'b10010100;
DRAM[51720] = 8'b10010100;
DRAM[51721] = 8'b10010100;
DRAM[51722] = 8'b10010101;
DRAM[51723] = 8'b10010101;
DRAM[51724] = 8'b10010101;
DRAM[51725] = 8'b10010101;
DRAM[51726] = 8'b10010110;
DRAM[51727] = 8'b10010110;
DRAM[51728] = 8'b10010010;
DRAM[51729] = 8'b10010011;
DRAM[51730] = 8'b10010100;
DRAM[51731] = 8'b10010101;
DRAM[51732] = 8'b10010111;
DRAM[51733] = 8'b10011011;
DRAM[51734] = 8'b10100001;
DRAM[51735] = 8'b10100110;
DRAM[51736] = 8'b10101011;
DRAM[51737] = 8'b10110110;
DRAM[51738] = 8'b11001001;
DRAM[51739] = 8'b11100000;
DRAM[51740] = 8'b11110100;
DRAM[51741] = 8'b11111110;
DRAM[51742] = 8'b11111110;
DRAM[51743] = 8'b11111010;
DRAM[51744] = 8'b11111101;
DRAM[51745] = 8'b11111101;
DRAM[51746] = 8'b11111101;
DRAM[51747] = 8'b11111101;
DRAM[51748] = 8'b11111011;
DRAM[51749] = 8'b11111010;
DRAM[51750] = 8'b11111000;
DRAM[51751] = 8'b11110111;
DRAM[51752] = 8'b11111000;
DRAM[51753] = 8'b11110110;
DRAM[51754] = 8'b11110100;
DRAM[51755] = 8'b11110010;
DRAM[51756] = 8'b11110000;
DRAM[51757] = 8'b11101101;
DRAM[51758] = 8'b11101000;
DRAM[51759] = 8'b11100100;
DRAM[51760] = 8'b11010100;
DRAM[51761] = 8'b11010001;
DRAM[51762] = 8'b11001110;
DRAM[51763] = 8'b11001101;
DRAM[51764] = 8'b11001100;
DRAM[51765] = 8'b11001010;
DRAM[51766] = 8'b11000111;
DRAM[51767] = 8'b11000101;
DRAM[51768] = 8'b11001001;
DRAM[51769] = 8'b11001100;
DRAM[51770] = 8'b11001101;
DRAM[51771] = 8'b11001001;
DRAM[51772] = 8'b11000110;
DRAM[51773] = 8'b11000111;
DRAM[51774] = 8'b11000110;
DRAM[51775] = 8'b11000100;
DRAM[51776] = 8'b11000001;
DRAM[51777] = 8'b10111001;
DRAM[51778] = 8'b10110110;
DRAM[51779] = 8'b10111100;
DRAM[51780] = 8'b11000011;
DRAM[51781] = 8'b11000001;
DRAM[51782] = 8'b10111011;
DRAM[51783] = 8'b10110110;
DRAM[51784] = 8'b11000000;
DRAM[51785] = 8'b10110111;
DRAM[51786] = 8'b10110010;
DRAM[51787] = 8'b10110100;
DRAM[51788] = 8'b10110110;
DRAM[51789] = 8'b10110101;
DRAM[51790] = 8'b10110010;
DRAM[51791] = 8'b10110000;
DRAM[51792] = 8'b10101011;
DRAM[51793] = 8'b10100111;
DRAM[51794] = 8'b10100010;
DRAM[51795] = 8'b10011101;
DRAM[51796] = 8'b10011000;
DRAM[51797] = 8'b10010010;
DRAM[51798] = 8'b10001011;
DRAM[51799] = 8'b10000110;
DRAM[51800] = 8'b10000110;
DRAM[51801] = 8'b10010010;
DRAM[51802] = 8'b10001000;
DRAM[51803] = 8'b10100010;
DRAM[51804] = 8'b10001101;
DRAM[51805] = 8'b10100000;
DRAM[51806] = 8'b10001010;
DRAM[51807] = 8'b10001101;
DRAM[51808] = 8'b10000010;
DRAM[51809] = 8'b10000000;
DRAM[51810] = 8'b10000010;
DRAM[51811] = 8'b1110101;
DRAM[51812] = 8'b1011001;
DRAM[51813] = 8'b1010100;
DRAM[51814] = 8'b1101001;
DRAM[51815] = 8'b1111010;
DRAM[51816] = 8'b1101110;
DRAM[51817] = 8'b1101000;
DRAM[51818] = 8'b1100111;
DRAM[51819] = 8'b1101100;
DRAM[51820] = 8'b1110000;
DRAM[51821] = 8'b1101101;
DRAM[51822] = 8'b1101000;
DRAM[51823] = 8'b1100101;
DRAM[51824] = 8'b1100011;
DRAM[51825] = 8'b1101000;
DRAM[51826] = 8'b1100001;
DRAM[51827] = 8'b1011011;
DRAM[51828] = 8'b1011110;
DRAM[51829] = 8'b1011100;
DRAM[51830] = 8'b1011011;
DRAM[51831] = 8'b1100011;
DRAM[51832] = 8'b1011101;
DRAM[51833] = 8'b1011101;
DRAM[51834] = 8'b1011110;
DRAM[51835] = 8'b1100001;
DRAM[51836] = 8'b1100100;
DRAM[51837] = 8'b1100010;
DRAM[51838] = 8'b1011011;
DRAM[51839] = 8'b1010101;
DRAM[51840] = 8'b1011111;
DRAM[51841] = 8'b1101011;
DRAM[51842] = 8'b1011101;
DRAM[51843] = 8'b1010110;
DRAM[51844] = 8'b1010011;
DRAM[51845] = 8'b1010100;
DRAM[51846] = 8'b1011101;
DRAM[51847] = 8'b1001111;
DRAM[51848] = 8'b1100010;
DRAM[51849] = 8'b1011011;
DRAM[51850] = 8'b1010111;
DRAM[51851] = 8'b1011010;
DRAM[51852] = 8'b1011111;
DRAM[51853] = 8'b1100011;
DRAM[51854] = 8'b1100110;
DRAM[51855] = 8'b1101010;
DRAM[51856] = 8'b1100110;
DRAM[51857] = 8'b1110110;
DRAM[51858] = 8'b1110111;
DRAM[51859] = 8'b1100110;
DRAM[51860] = 8'b1100011;
DRAM[51861] = 8'b1110010;
DRAM[51862] = 8'b1111000;
DRAM[51863] = 8'b1110000;
DRAM[51864] = 8'b1101001;
DRAM[51865] = 8'b1101101;
DRAM[51866] = 8'b1110000;
DRAM[51867] = 8'b1110000;
DRAM[51868] = 8'b1110011;
DRAM[51869] = 8'b1111000;
DRAM[51870] = 8'b1111011;
DRAM[51871] = 8'b1111011;
DRAM[51872] = 8'b10000010;
DRAM[51873] = 8'b10000001;
DRAM[51874] = 8'b10000011;
DRAM[51875] = 8'b10001011;
DRAM[51876] = 8'b10010100;
DRAM[51877] = 8'b10010110;
DRAM[51878] = 8'b10010001;
DRAM[51879] = 8'b10001010;
DRAM[51880] = 8'b10010011;
DRAM[51881] = 8'b10010010;
DRAM[51882] = 8'b10010001;
DRAM[51883] = 8'b10010100;
DRAM[51884] = 8'b10011010;
DRAM[51885] = 8'b10100000;
DRAM[51886] = 8'b10100011;
DRAM[51887] = 8'b10100101;
DRAM[51888] = 8'b10100101;
DRAM[51889] = 8'b10100110;
DRAM[51890] = 8'b10101100;
DRAM[51891] = 8'b10110100;
DRAM[51892] = 8'b10111010;
DRAM[51893] = 8'b10111100;
DRAM[51894] = 8'b11000011;
DRAM[51895] = 8'b11001010;
DRAM[51896] = 8'b11011111;
DRAM[51897] = 8'b11100011;
DRAM[51898] = 8'b11100110;
DRAM[51899] = 8'b11100111;
DRAM[51900] = 8'b11100101;
DRAM[51901] = 8'b11100110;
DRAM[51902] = 8'b11101001;
DRAM[51903] = 8'b11101101;
DRAM[51904] = 8'b11111100;
DRAM[51905] = 8'b11111000;
DRAM[51906] = 8'b11110001;
DRAM[51907] = 8'b11100111;
DRAM[51908] = 8'b11011010;
DRAM[51909] = 8'b11001010;
DRAM[51910] = 8'b10111010;
DRAM[51911] = 8'b10110001;
DRAM[51912] = 8'b10100001;
DRAM[51913] = 8'b10011000;
DRAM[51914] = 8'b10001111;
DRAM[51915] = 8'b10001101;
DRAM[51916] = 8'b10001001;
DRAM[51917] = 8'b10000010;
DRAM[51918] = 8'b1111101;
DRAM[51919] = 8'b1111011;
DRAM[51920] = 8'b1111100;
DRAM[51921] = 8'b1111001;
DRAM[51922] = 8'b1110101;
DRAM[51923] = 8'b1110011;
DRAM[51924] = 8'b1110010;
DRAM[51925] = 8'b1110000;
DRAM[51926] = 8'b1101110;
DRAM[51927] = 8'b1101100;
DRAM[51928] = 8'b1101111;
DRAM[51929] = 8'b1101101;
DRAM[51930] = 8'b1101101;
DRAM[51931] = 8'b1101110;
DRAM[51932] = 8'b1110001;
DRAM[51933] = 8'b1110010;
DRAM[51934] = 8'b1110010;
DRAM[51935] = 8'b1110000;
DRAM[51936] = 8'b1110000;
DRAM[51937] = 8'b1110001;
DRAM[51938] = 8'b1110010;
DRAM[51939] = 8'b1110100;
DRAM[51940] = 8'b1110110;
DRAM[51941] = 8'b1111000;
DRAM[51942] = 8'b1111001;
DRAM[51943] = 8'b1111010;
DRAM[51944] = 8'b1111000;
DRAM[51945] = 8'b1111000;
DRAM[51946] = 8'b1111000;
DRAM[51947] = 8'b1111000;
DRAM[51948] = 8'b1111000;
DRAM[51949] = 8'b1111000;
DRAM[51950] = 8'b1111000;
DRAM[51951] = 8'b1111000;
DRAM[51952] = 8'b1110110;
DRAM[51953] = 8'b1110101;
DRAM[51954] = 8'b1110101;
DRAM[51955] = 8'b1110100;
DRAM[51956] = 8'b1110011;
DRAM[51957] = 8'b1110010;
DRAM[51958] = 8'b1110010;
DRAM[51959] = 8'b1110001;
DRAM[51960] = 8'b1110100;
DRAM[51961] = 8'b1110011;
DRAM[51962] = 8'b1110011;
DRAM[51963] = 8'b1110011;
DRAM[51964] = 8'b1110011;
DRAM[51965] = 8'b1110100;
DRAM[51966] = 8'b1110101;
DRAM[51967] = 8'b1110110;
DRAM[51968] = 8'b10001100;
DRAM[51969] = 8'b10001100;
DRAM[51970] = 8'b10001101;
DRAM[51971] = 8'b10001110;
DRAM[51972] = 8'b10010000;
DRAM[51973] = 8'b10010010;
DRAM[51974] = 8'b10010011;
DRAM[51975] = 8'b10010100;
DRAM[51976] = 8'b10010101;
DRAM[51977] = 8'b10010101;
DRAM[51978] = 8'b10010101;
DRAM[51979] = 8'b10010101;
DRAM[51980] = 8'b10010101;
DRAM[51981] = 8'b10010101;
DRAM[51982] = 8'b10010101;
DRAM[51983] = 8'b10010101;
DRAM[51984] = 8'b10010011;
DRAM[51985] = 8'b10010100;
DRAM[51986] = 8'b10010101;
DRAM[51987] = 8'b10010101;
DRAM[51988] = 8'b10010111;
DRAM[51989] = 8'b10011011;
DRAM[51990] = 8'b10100001;
DRAM[51991] = 8'b10100110;
DRAM[51992] = 8'b10100110;
DRAM[51993] = 8'b10111001;
DRAM[51994] = 8'b11010010;
DRAM[51995] = 8'b11101000;
DRAM[51996] = 8'b11110111;
DRAM[51997] = 8'b11111111;
DRAM[51998] = 8'b11111111;
DRAM[51999] = 8'b11111011;
DRAM[52000] = 8'b11111101;
DRAM[52001] = 8'b11111101;
DRAM[52002] = 8'b11111100;
DRAM[52003] = 8'b11111100;
DRAM[52004] = 8'b11111011;
DRAM[52005] = 8'b11111010;
DRAM[52006] = 8'b11111001;
DRAM[52007] = 8'b11111001;
DRAM[52008] = 8'b11111000;
DRAM[52009] = 8'b11110110;
DRAM[52010] = 8'b11110100;
DRAM[52011] = 8'b11110011;
DRAM[52012] = 8'b11110001;
DRAM[52013] = 8'b11101101;
DRAM[52014] = 8'b11101001;
DRAM[52015] = 8'b11100101;
DRAM[52016] = 8'b11101000;
DRAM[52017] = 8'b11100101;
DRAM[52018] = 8'b11011111;
DRAM[52019] = 8'b11011010;
DRAM[52020] = 8'b11010110;
DRAM[52021] = 8'b11010000;
DRAM[52022] = 8'b11001010;
DRAM[52023] = 8'b11000110;
DRAM[52024] = 8'b11001000;
DRAM[52025] = 8'b11001001;
DRAM[52026] = 8'b11001010;
DRAM[52027] = 8'b11001011;
DRAM[52028] = 8'b11001101;
DRAM[52029] = 8'b11001100;
DRAM[52030] = 8'b11000111;
DRAM[52031] = 8'b11000001;
DRAM[52032] = 8'b11000010;
DRAM[52033] = 8'b10111000;
DRAM[52034] = 8'b10110010;
DRAM[52035] = 8'b10111000;
DRAM[52036] = 8'b11000010;
DRAM[52037] = 8'b11000111;
DRAM[52038] = 8'b11000111;
DRAM[52039] = 8'b11000111;
DRAM[52040] = 8'b11000001;
DRAM[52041] = 8'b10101110;
DRAM[52042] = 8'b10100011;
DRAM[52043] = 8'b10101100;
DRAM[52044] = 8'b10111000;
DRAM[52045] = 8'b10110110;
DRAM[52046] = 8'b10101111;
DRAM[52047] = 8'b10101011;
DRAM[52048] = 8'b10101000;
DRAM[52049] = 8'b10100010;
DRAM[52050] = 8'b10011001;
DRAM[52051] = 8'b10010001;
DRAM[52052] = 8'b10001011;
DRAM[52053] = 8'b10000101;
DRAM[52054] = 8'b10000001;
DRAM[52055] = 8'b1111110;
DRAM[52056] = 8'b1111110;
DRAM[52057] = 8'b10001010;
DRAM[52058] = 8'b10001100;
DRAM[52059] = 8'b10011010;
DRAM[52060] = 8'b10010000;
DRAM[52061] = 8'b10011001;
DRAM[52062] = 8'b10001100;
DRAM[52063] = 8'b10001011;
DRAM[52064] = 8'b10001100;
DRAM[52065] = 8'b10000100;
DRAM[52066] = 8'b1111111;
DRAM[52067] = 8'b1101101;
DRAM[52068] = 8'b1010101;
DRAM[52069] = 8'b1010110;
DRAM[52070] = 8'b1101100;
DRAM[52071] = 8'b1111011;
DRAM[52072] = 8'b1110111;
DRAM[52073] = 8'b1101011;
DRAM[52074] = 8'b1100111;
DRAM[52075] = 8'b1101111;
DRAM[52076] = 8'b1110010;
DRAM[52077] = 8'b1101010;
DRAM[52078] = 8'b1100010;
DRAM[52079] = 8'b1100000;
DRAM[52080] = 8'b1011111;
DRAM[52081] = 8'b1101001;
DRAM[52082] = 8'b1100010;
DRAM[52083] = 8'b1011000;
DRAM[52084] = 8'b1011101;
DRAM[52085] = 8'b1100001;
DRAM[52086] = 8'b1011111;
DRAM[52087] = 8'b1100000;
DRAM[52088] = 8'b1011111;
DRAM[52089] = 8'b1011111;
DRAM[52090] = 8'b1100001;
DRAM[52091] = 8'b1100100;
DRAM[52092] = 8'b1100110;
DRAM[52093] = 8'b1100010;
DRAM[52094] = 8'b1011001;
DRAM[52095] = 8'b1010010;
DRAM[52096] = 8'b1011110;
DRAM[52097] = 8'b1101000;
DRAM[52098] = 8'b1011011;
DRAM[52099] = 8'b1010110;
DRAM[52100] = 8'b1010100;
DRAM[52101] = 8'b1010101;
DRAM[52102] = 8'b1011111;
DRAM[52103] = 8'b1010011;
DRAM[52104] = 8'b1100011;
DRAM[52105] = 8'b1011001;
DRAM[52106] = 8'b1010010;
DRAM[52107] = 8'b1010100;
DRAM[52108] = 8'b1011010;
DRAM[52109] = 8'b1011110;
DRAM[52110] = 8'b1100000;
DRAM[52111] = 8'b1100011;
DRAM[52112] = 8'b1011110;
DRAM[52113] = 8'b1101011;
DRAM[52114] = 8'b1101111;
DRAM[52115] = 8'b1100100;
DRAM[52116] = 8'b1011110;
DRAM[52117] = 8'b1100101;
DRAM[52118] = 8'b1101110;
DRAM[52119] = 8'b1110000;
DRAM[52120] = 8'b1100101;
DRAM[52121] = 8'b1101110;
DRAM[52122] = 8'b1110100;
DRAM[52123] = 8'b1110010;
DRAM[52124] = 8'b1110010;
DRAM[52125] = 8'b1111000;
DRAM[52126] = 8'b1111100;
DRAM[52127] = 8'b1111100;
DRAM[52128] = 8'b10000011;
DRAM[52129] = 8'b10001000;
DRAM[52130] = 8'b10001010;
DRAM[52131] = 8'b10001011;
DRAM[52132] = 8'b10010010;
DRAM[52133] = 8'b10011011;
DRAM[52134] = 8'b10011011;
DRAM[52135] = 8'b10010011;
DRAM[52136] = 8'b10010100;
DRAM[52137] = 8'b10010101;
DRAM[52138] = 8'b10010111;
DRAM[52139] = 8'b10011000;
DRAM[52140] = 8'b10011010;
DRAM[52141] = 8'b10100000;
DRAM[52142] = 8'b10101000;
DRAM[52143] = 8'b10101101;
DRAM[52144] = 8'b10110001;
DRAM[52145] = 8'b10110001;
DRAM[52146] = 8'b10110110;
DRAM[52147] = 8'b10111101;
DRAM[52148] = 8'b10111111;
DRAM[52149] = 8'b10111110;
DRAM[52150] = 8'b11000000;
DRAM[52151] = 8'b11000101;
DRAM[52152] = 8'b11001100;
DRAM[52153] = 8'b11010011;
DRAM[52154] = 8'b11011111;
DRAM[52155] = 8'b11101000;
DRAM[52156] = 8'b11101101;
DRAM[52157] = 8'b11101101;
DRAM[52158] = 8'b11101011;
DRAM[52159] = 8'b11101001;
DRAM[52160] = 8'b11101100;
DRAM[52161] = 8'b11101100;
DRAM[52162] = 8'b11101100;
DRAM[52163] = 8'b11101000;
DRAM[52164] = 8'b11011101;
DRAM[52165] = 8'b11001010;
DRAM[52166] = 8'b10110101;
DRAM[52167] = 8'b10100111;
DRAM[52168] = 8'b10011111;
DRAM[52169] = 8'b10010110;
DRAM[52170] = 8'b10001101;
DRAM[52171] = 8'b10001010;
DRAM[52172] = 8'b10000111;
DRAM[52173] = 8'b10000001;
DRAM[52174] = 8'b1111100;
DRAM[52175] = 8'b1111011;
DRAM[52176] = 8'b1111001;
DRAM[52177] = 8'b1110111;
DRAM[52178] = 8'b1110011;
DRAM[52179] = 8'b1110001;
DRAM[52180] = 8'b1110001;
DRAM[52181] = 8'b1110000;
DRAM[52182] = 8'b1101110;
DRAM[52183] = 8'b1101100;
DRAM[52184] = 8'b1101110;
DRAM[52185] = 8'b1101101;
DRAM[52186] = 8'b1101100;
DRAM[52187] = 8'b1101101;
DRAM[52188] = 8'b1110000;
DRAM[52189] = 8'b1110001;
DRAM[52190] = 8'b1110001;
DRAM[52191] = 8'b1110000;
DRAM[52192] = 8'b1110000;
DRAM[52193] = 8'b1110001;
DRAM[52194] = 8'b1110010;
DRAM[52195] = 8'b1110100;
DRAM[52196] = 8'b1110110;
DRAM[52197] = 8'b1111000;
DRAM[52198] = 8'b1111001;
DRAM[52199] = 8'b1111010;
DRAM[52200] = 8'b1111000;
DRAM[52201] = 8'b1111000;
DRAM[52202] = 8'b1111000;
DRAM[52203] = 8'b1111000;
DRAM[52204] = 8'b1110111;
DRAM[52205] = 8'b1110111;
DRAM[52206] = 8'b1110111;
DRAM[52207] = 8'b1110111;
DRAM[52208] = 8'b1110101;
DRAM[52209] = 8'b1110101;
DRAM[52210] = 8'b1110100;
DRAM[52211] = 8'b1110011;
DRAM[52212] = 8'b1110011;
DRAM[52213] = 8'b1110010;
DRAM[52214] = 8'b1110001;
DRAM[52215] = 8'b1110001;
DRAM[52216] = 8'b1110010;
DRAM[52217] = 8'b1110010;
DRAM[52218] = 8'b1110010;
DRAM[52219] = 8'b1110010;
DRAM[52220] = 8'b1110011;
DRAM[52221] = 8'b1110011;
DRAM[52222] = 8'b1110100;
DRAM[52223] = 8'b1110100;
DRAM[52224] = 8'b10001100;
DRAM[52225] = 8'b10001101;
DRAM[52226] = 8'b10001110;
DRAM[52227] = 8'b10010000;
DRAM[52228] = 8'b10010010;
DRAM[52229] = 8'b10010011;
DRAM[52230] = 8'b10010100;
DRAM[52231] = 8'b10010100;
DRAM[52232] = 8'b10010101;
DRAM[52233] = 8'b10010101;
DRAM[52234] = 8'b10010101;
DRAM[52235] = 8'b10010101;
DRAM[52236] = 8'b10010101;
DRAM[52237] = 8'b10010101;
DRAM[52238] = 8'b10010101;
DRAM[52239] = 8'b10010101;
DRAM[52240] = 8'b10010100;
DRAM[52241] = 8'b10010101;
DRAM[52242] = 8'b10010101;
DRAM[52243] = 8'b10010101;
DRAM[52244] = 8'b10010110;
DRAM[52245] = 8'b10011010;
DRAM[52246] = 8'b10011111;
DRAM[52247] = 8'b10100011;
DRAM[52248] = 8'b10101011;
DRAM[52249] = 8'b11000011;
DRAM[52250] = 8'b11100000;
DRAM[52251] = 8'b11110001;
DRAM[52252] = 8'b11111011;
DRAM[52253] = 8'b11111111;
DRAM[52254] = 8'b11111111;
DRAM[52255] = 8'b11111011;
DRAM[52256] = 8'b11111100;
DRAM[52257] = 8'b11111100;
DRAM[52258] = 8'b11111100;
DRAM[52259] = 8'b11111011;
DRAM[52260] = 8'b11111011;
DRAM[52261] = 8'b11111011;
DRAM[52262] = 8'b11111011;
DRAM[52263] = 8'b11111011;
DRAM[52264] = 8'b11111001;
DRAM[52265] = 8'b11110111;
DRAM[52266] = 8'b11110101;
DRAM[52267] = 8'b11110100;
DRAM[52268] = 8'b11110011;
DRAM[52269] = 8'b11110000;
DRAM[52270] = 8'b11101011;
DRAM[52271] = 8'b11101000;
DRAM[52272] = 8'b11101110;
DRAM[52273] = 8'b11101011;
DRAM[52274] = 8'b11101000;
DRAM[52275] = 8'b11100101;
DRAM[52276] = 8'b11100001;
DRAM[52277] = 8'b11011101;
DRAM[52278] = 8'b11011000;
DRAM[52279] = 8'b11010100;
DRAM[52280] = 8'b11000111;
DRAM[52281] = 8'b11000100;
DRAM[52282] = 8'b11000100;
DRAM[52283] = 8'b11001011;
DRAM[52284] = 8'b11010010;
DRAM[52285] = 8'b11010000;
DRAM[52286] = 8'b11000101;
DRAM[52287] = 8'b10111100;
DRAM[52288] = 8'b10111111;
DRAM[52289] = 8'b10111100;
DRAM[52290] = 8'b10111101;
DRAM[52291] = 8'b11000011;
DRAM[52292] = 8'b11000100;
DRAM[52293] = 8'b10111101;
DRAM[52294] = 8'b10110110;
DRAM[52295] = 8'b10110011;
DRAM[52296] = 8'b10101111;
DRAM[52297] = 8'b10101010;
DRAM[52298] = 8'b10101010;
DRAM[52299] = 8'b10101101;
DRAM[52300] = 8'b10101000;
DRAM[52301] = 8'b10011110;
DRAM[52302] = 8'b10011110;
DRAM[52303] = 8'b10100110;
DRAM[52304] = 8'b10100110;
DRAM[52305] = 8'b10011111;
DRAM[52306] = 8'b10010101;
DRAM[52307] = 8'b10001100;
DRAM[52308] = 8'b10001000;
DRAM[52309] = 8'b10000110;
DRAM[52310] = 8'b10000110;
DRAM[52311] = 8'b10000110;
DRAM[52312] = 8'b1111101;
DRAM[52313] = 8'b10000111;
DRAM[52314] = 8'b10011011;
DRAM[52315] = 8'b10010000;
DRAM[52316] = 8'b10011000;
DRAM[52317] = 8'b10001100;
DRAM[52318] = 8'b10010010;
DRAM[52319] = 8'b10001011;
DRAM[52320] = 8'b10010000;
DRAM[52321] = 8'b10000001;
DRAM[52322] = 8'b1110100;
DRAM[52323] = 8'b1100100;
DRAM[52324] = 8'b1010110;
DRAM[52325] = 8'b1011110;
DRAM[52326] = 8'b1110001;
DRAM[52327] = 8'b1110111;
DRAM[52328] = 8'b1111010;
DRAM[52329] = 8'b1101110;
DRAM[52330] = 8'b1101001;
DRAM[52331] = 8'b1110000;
DRAM[52332] = 8'b1110010;
DRAM[52333] = 8'b1101001;
DRAM[52334] = 8'b1100000;
DRAM[52335] = 8'b1011110;
DRAM[52336] = 8'b1011110;
DRAM[52337] = 8'b1101001;
DRAM[52338] = 8'b1100010;
DRAM[52339] = 8'b1010111;
DRAM[52340] = 8'b1011101;
DRAM[52341] = 8'b1100011;
DRAM[52342] = 8'b1100000;
DRAM[52343] = 8'b1011110;
DRAM[52344] = 8'b1100011;
DRAM[52345] = 8'b1100011;
DRAM[52346] = 8'b1100100;
DRAM[52347] = 8'b1100110;
DRAM[52348] = 8'b1100110;
DRAM[52349] = 8'b1100000;
DRAM[52350] = 8'b1010110;
DRAM[52351] = 8'b1001110;
DRAM[52352] = 8'b1011100;
DRAM[52353] = 8'b1100100;
DRAM[52354] = 8'b1010111;
DRAM[52355] = 8'b1010101;
DRAM[52356] = 8'b1010100;
DRAM[52357] = 8'b1010101;
DRAM[52358] = 8'b1100000;
DRAM[52359] = 8'b1010111;
DRAM[52360] = 8'b1100101;
DRAM[52361] = 8'b1011010;
DRAM[52362] = 8'b1010010;
DRAM[52363] = 8'b1010100;
DRAM[52364] = 8'b1011000;
DRAM[52365] = 8'b1011010;
DRAM[52366] = 8'b1011011;
DRAM[52367] = 8'b1011101;
DRAM[52368] = 8'b1100110;
DRAM[52369] = 8'b1100110;
DRAM[52370] = 8'b1101101;
DRAM[52371] = 8'b1110011;
DRAM[52372] = 8'b1101101;
DRAM[52373] = 8'b1100101;
DRAM[52374] = 8'b1101100;
DRAM[52375] = 8'b1111011;
DRAM[52376] = 8'b1101001;
DRAM[52377] = 8'b1101111;
DRAM[52378] = 8'b1110011;
DRAM[52379] = 8'b1110010;
DRAM[52380] = 8'b1110010;
DRAM[52381] = 8'b1110111;
DRAM[52382] = 8'b1111100;
DRAM[52383] = 8'b1111110;
DRAM[52384] = 8'b1111101;
DRAM[52385] = 8'b10001001;
DRAM[52386] = 8'b10001110;
DRAM[52387] = 8'b10001010;
DRAM[52388] = 8'b10001100;
DRAM[52389] = 8'b10011000;
DRAM[52390] = 8'b10011101;
DRAM[52391] = 8'b10011010;
DRAM[52392] = 8'b10011010;
DRAM[52393] = 8'b10011101;
DRAM[52394] = 8'b10011111;
DRAM[52395] = 8'b10011111;
DRAM[52396] = 8'b10011101;
DRAM[52397] = 8'b10100000;
DRAM[52398] = 8'b10101000;
DRAM[52399] = 8'b10101110;
DRAM[52400] = 8'b10110100;
DRAM[52401] = 8'b10110110;
DRAM[52402] = 8'b10111011;
DRAM[52403] = 8'b11000011;
DRAM[52404] = 8'b11000110;
DRAM[52405] = 8'b11000101;
DRAM[52406] = 8'b11000111;
DRAM[52407] = 8'b11001100;
DRAM[52408] = 8'b11000011;
DRAM[52409] = 8'b11001001;
DRAM[52410] = 8'b11010011;
DRAM[52411] = 8'b11011111;
DRAM[52412] = 8'b11101000;
DRAM[52413] = 8'b11101100;
DRAM[52414] = 8'b11101011;
DRAM[52415] = 8'b11101001;
DRAM[52416] = 8'b11101110;
DRAM[52417] = 8'b11101101;
DRAM[52418] = 8'b11101011;
DRAM[52419] = 8'b11100011;
DRAM[52420] = 8'b11010101;
DRAM[52421] = 8'b11000010;
DRAM[52422] = 8'b10101110;
DRAM[52423] = 8'b10100001;
DRAM[52424] = 8'b10100000;
DRAM[52425] = 8'b10010100;
DRAM[52426] = 8'b10001001;
DRAM[52427] = 8'b10000100;
DRAM[52428] = 8'b10000001;
DRAM[52429] = 8'b1111101;
DRAM[52430] = 8'b1111011;
DRAM[52431] = 8'b1111100;
DRAM[52432] = 8'b1110110;
DRAM[52433] = 8'b1110100;
DRAM[52434] = 8'b1110001;
DRAM[52435] = 8'b1110001;
DRAM[52436] = 8'b1110001;
DRAM[52437] = 8'b1110001;
DRAM[52438] = 8'b1110000;
DRAM[52439] = 8'b1101111;
DRAM[52440] = 8'b1101111;
DRAM[52441] = 8'b1101101;
DRAM[52442] = 8'b1101100;
DRAM[52443] = 8'b1101101;
DRAM[52444] = 8'b1101111;
DRAM[52445] = 8'b1110001;
DRAM[52446] = 8'b1110001;
DRAM[52447] = 8'b1110001;
DRAM[52448] = 8'b1110001;
DRAM[52449] = 8'b1110001;
DRAM[52450] = 8'b1110010;
DRAM[52451] = 8'b1110100;
DRAM[52452] = 8'b1110110;
DRAM[52453] = 8'b1111000;
DRAM[52454] = 8'b1111001;
DRAM[52455] = 8'b1111001;
DRAM[52456] = 8'b1111000;
DRAM[52457] = 8'b1111000;
DRAM[52458] = 8'b1110111;
DRAM[52459] = 8'b1110111;
DRAM[52460] = 8'b1110110;
DRAM[52461] = 8'b1110110;
DRAM[52462] = 8'b1110101;
DRAM[52463] = 8'b1110101;
DRAM[52464] = 8'b1110101;
DRAM[52465] = 8'b1110101;
DRAM[52466] = 8'b1110100;
DRAM[52467] = 8'b1110011;
DRAM[52468] = 8'b1110011;
DRAM[52469] = 8'b1110010;
DRAM[52470] = 8'b1110001;
DRAM[52471] = 8'b1110001;
DRAM[52472] = 8'b1110000;
DRAM[52473] = 8'b1110000;
DRAM[52474] = 8'b1110001;
DRAM[52475] = 8'b1110001;
DRAM[52476] = 8'b1110010;
DRAM[52477] = 8'b1110010;
DRAM[52478] = 8'b1110010;
DRAM[52479] = 8'b1110010;
DRAM[52480] = 8'b10001100;
DRAM[52481] = 8'b10001101;
DRAM[52482] = 8'b10001111;
DRAM[52483] = 8'b10010001;
DRAM[52484] = 8'b10010011;
DRAM[52485] = 8'b10010100;
DRAM[52486] = 8'b10010100;
DRAM[52487] = 8'b10010100;
DRAM[52488] = 8'b10010110;
DRAM[52489] = 8'b10010110;
DRAM[52490] = 8'b10010101;
DRAM[52491] = 8'b10010101;
DRAM[52492] = 8'b10010101;
DRAM[52493] = 8'b10010101;
DRAM[52494] = 8'b10010100;
DRAM[52495] = 8'b10010100;
DRAM[52496] = 8'b10010101;
DRAM[52497] = 8'b10010110;
DRAM[52498] = 8'b10010110;
DRAM[52499] = 8'b10010101;
DRAM[52500] = 8'b10010110;
DRAM[52501] = 8'b10011010;
DRAM[52502] = 8'b10011111;
DRAM[52503] = 8'b10100011;
DRAM[52504] = 8'b10111000;
DRAM[52505] = 8'b11010100;
DRAM[52506] = 8'b11110001;
DRAM[52507] = 8'b11111100;
DRAM[52508] = 8'b11111101;
DRAM[52509] = 8'b11111111;
DRAM[52510] = 8'b11111110;
DRAM[52511] = 8'b11111100;
DRAM[52512] = 8'b11111101;
DRAM[52513] = 8'b11111100;
DRAM[52514] = 8'b11111011;
DRAM[52515] = 8'b11111001;
DRAM[52516] = 8'b11111001;
DRAM[52517] = 8'b11111000;
DRAM[52518] = 8'b11111001;
DRAM[52519] = 8'b11111001;
DRAM[52520] = 8'b11110111;
DRAM[52521] = 8'b11110110;
DRAM[52522] = 8'b11110101;
DRAM[52523] = 8'b11110100;
DRAM[52524] = 8'b11110100;
DRAM[52525] = 8'b11110001;
DRAM[52526] = 8'b11101101;
DRAM[52527] = 8'b11101010;
DRAM[52528] = 8'b11100110;
DRAM[52529] = 8'b11100011;
DRAM[52530] = 8'b11100000;
DRAM[52531] = 8'b11011110;
DRAM[52532] = 8'b11011010;
DRAM[52533] = 8'b11010101;
DRAM[52534] = 8'b11010000;
DRAM[52535] = 8'b11001011;
DRAM[52536] = 8'b11001001;
DRAM[52537] = 8'b11000011;
DRAM[52538] = 8'b11000010;
DRAM[52539] = 8'b11001010;
DRAM[52540] = 8'b11010000;
DRAM[52541] = 8'b11001100;
DRAM[52542] = 8'b11000001;
DRAM[52543] = 8'b10111010;
DRAM[52544] = 8'b11000111;
DRAM[52545] = 8'b11000100;
DRAM[52546] = 8'b11000011;
DRAM[52547] = 8'b11000010;
DRAM[52548] = 8'b10111101;
DRAM[52549] = 8'b10110100;
DRAM[52550] = 8'b10110001;
DRAM[52551] = 8'b10110010;
DRAM[52552] = 8'b10101010;
DRAM[52553] = 8'b10100111;
DRAM[52554] = 8'b10100111;
DRAM[52555] = 8'b10101001;
DRAM[52556] = 8'b10101001;
DRAM[52557] = 8'b10100100;
DRAM[52558] = 8'b10100001;
DRAM[52559] = 8'b10100001;
DRAM[52560] = 8'b10011111;
DRAM[52561] = 8'b10011010;
DRAM[52562] = 8'b10010010;
DRAM[52563] = 8'b10001101;
DRAM[52564] = 8'b10001100;
DRAM[52565] = 8'b10001101;
DRAM[52566] = 8'b10001111;
DRAM[52567] = 8'b10010000;
DRAM[52568] = 8'b10000101;
DRAM[52569] = 8'b10001100;
DRAM[52570] = 8'b10100101;
DRAM[52571] = 8'b10001011;
DRAM[52572] = 8'b10011010;
DRAM[52573] = 8'b10000100;
DRAM[52574] = 8'b10010100;
DRAM[52575] = 8'b10001001;
DRAM[52576] = 8'b10000111;
DRAM[52577] = 8'b1110100;
DRAM[52578] = 8'b1100101;
DRAM[52579] = 8'b1011010;
DRAM[52580] = 8'b1010111;
DRAM[52581] = 8'b1100111;
DRAM[52582] = 8'b1110111;
DRAM[52583] = 8'b1110101;
DRAM[52584] = 8'b1110101;
DRAM[52585] = 8'b1101111;
DRAM[52586] = 8'b1101100;
DRAM[52587] = 8'b1101111;
DRAM[52588] = 8'b1110000;
DRAM[52589] = 8'b1101011;
DRAM[52590] = 8'b1100100;
DRAM[52591] = 8'b1100000;
DRAM[52592] = 8'b1100001;
DRAM[52593] = 8'b1101001;
DRAM[52594] = 8'b1100010;
DRAM[52595] = 8'b1011010;
DRAM[52596] = 8'b1100000;
DRAM[52597] = 8'b1100100;
DRAM[52598] = 8'b1100000;
DRAM[52599] = 8'b1011111;
DRAM[52600] = 8'b1100110;
DRAM[52601] = 8'b1100101;
DRAM[52602] = 8'b1100101;
DRAM[52603] = 8'b1100110;
DRAM[52604] = 8'b1100101;
DRAM[52605] = 8'b1011110;
DRAM[52606] = 8'b1010100;
DRAM[52607] = 8'b1001011;
DRAM[52608] = 8'b1011011;
DRAM[52609] = 8'b1100001;
DRAM[52610] = 8'b1010100;
DRAM[52611] = 8'b1010011;
DRAM[52612] = 8'b1010010;
DRAM[52613] = 8'b1010010;
DRAM[52614] = 8'b1011110;
DRAM[52615] = 8'b1010111;
DRAM[52616] = 8'b1100101;
DRAM[52617] = 8'b1011110;
DRAM[52618] = 8'b1011001;
DRAM[52619] = 8'b1011011;
DRAM[52620] = 8'b1011101;
DRAM[52621] = 8'b1011100;
DRAM[52622] = 8'b1011100;
DRAM[52623] = 8'b1011110;
DRAM[52624] = 8'b1101001;
DRAM[52625] = 8'b1100001;
DRAM[52626] = 8'b1100111;
DRAM[52627] = 8'b1110111;
DRAM[52628] = 8'b1110110;
DRAM[52629] = 8'b1100111;
DRAM[52630] = 8'b1101011;
DRAM[52631] = 8'b1111101;
DRAM[52632] = 8'b1101101;
DRAM[52633] = 8'b1101100;
DRAM[52634] = 8'b1101110;
DRAM[52635] = 8'b1110011;
DRAM[52636] = 8'b1110101;
DRAM[52637] = 8'b1110110;
DRAM[52638] = 8'b1111011;
DRAM[52639] = 8'b10000001;
DRAM[52640] = 8'b1111101;
DRAM[52641] = 8'b10001001;
DRAM[52642] = 8'b10010000;
DRAM[52643] = 8'b10001101;
DRAM[52644] = 8'b10001110;
DRAM[52645] = 8'b10010111;
DRAM[52646] = 8'b10100000;
DRAM[52647] = 8'b10100010;
DRAM[52648] = 8'b10100010;
DRAM[52649] = 8'b10100110;
DRAM[52650] = 8'b10101001;
DRAM[52651] = 8'b10100111;
DRAM[52652] = 8'b10100011;
DRAM[52653] = 8'b10100010;
DRAM[52654] = 8'b10100101;
DRAM[52655] = 8'b10101010;
DRAM[52656] = 8'b10101111;
DRAM[52657] = 8'b10110001;
DRAM[52658] = 8'b10111001;
DRAM[52659] = 8'b11000100;
DRAM[52660] = 8'b11001010;
DRAM[52661] = 8'b11001101;
DRAM[52662] = 8'b11010010;
DRAM[52663] = 8'b11011001;
DRAM[52664] = 8'b11001111;
DRAM[52665] = 8'b11001101;
DRAM[52666] = 8'b11001100;
DRAM[52667] = 8'b11010010;
DRAM[52668] = 8'b11011011;
DRAM[52669] = 8'b11100101;
DRAM[52670] = 8'b11101010;
DRAM[52671] = 8'b11101100;
DRAM[52672] = 8'b11110010;
DRAM[52673] = 8'b11101110;
DRAM[52674] = 8'b11100101;
DRAM[52675] = 8'b11011000;
DRAM[52676] = 8'b11001001;
DRAM[52677] = 8'b10111100;
DRAM[52678] = 8'b10110100;
DRAM[52679] = 8'b10110000;
DRAM[52680] = 8'b10100000;
DRAM[52681] = 8'b10010011;
DRAM[52682] = 8'b10000110;
DRAM[52683] = 8'b1111111;
DRAM[52684] = 8'b1111101;
DRAM[52685] = 8'b1111010;
DRAM[52686] = 8'b1111011;
DRAM[52687] = 8'b1111110;
DRAM[52688] = 8'b1110110;
DRAM[52689] = 8'b1110100;
DRAM[52690] = 8'b1110010;
DRAM[52691] = 8'b1110010;
DRAM[52692] = 8'b1110011;
DRAM[52693] = 8'b1110011;
DRAM[52694] = 8'b1110011;
DRAM[52695] = 8'b1110010;
DRAM[52696] = 8'b1110000;
DRAM[52697] = 8'b1101110;
DRAM[52698] = 8'b1101100;
DRAM[52699] = 8'b1101101;
DRAM[52700] = 8'b1101111;
DRAM[52701] = 8'b1110001;
DRAM[52702] = 8'b1110010;
DRAM[52703] = 8'b1110010;
DRAM[52704] = 8'b1110010;
DRAM[52705] = 8'b1110011;
DRAM[52706] = 8'b1110011;
DRAM[52707] = 8'b1110100;
DRAM[52708] = 8'b1110110;
DRAM[52709] = 8'b1110111;
DRAM[52710] = 8'b1110111;
DRAM[52711] = 8'b1111000;
DRAM[52712] = 8'b1111000;
DRAM[52713] = 8'b1110111;
DRAM[52714] = 8'b1110111;
DRAM[52715] = 8'b1110110;
DRAM[52716] = 8'b1110101;
DRAM[52717] = 8'b1110101;
DRAM[52718] = 8'b1110100;
DRAM[52719] = 8'b1110100;
DRAM[52720] = 8'b1110101;
DRAM[52721] = 8'b1110100;
DRAM[52722] = 8'b1110100;
DRAM[52723] = 8'b1110011;
DRAM[52724] = 8'b1110010;
DRAM[52725] = 8'b1110001;
DRAM[52726] = 8'b1110001;
DRAM[52727] = 8'b1110000;
DRAM[52728] = 8'b1101110;
DRAM[52729] = 8'b1101111;
DRAM[52730] = 8'b1110000;
DRAM[52731] = 8'b1110001;
DRAM[52732] = 8'b1110001;
DRAM[52733] = 8'b1110001;
DRAM[52734] = 8'b1110001;
DRAM[52735] = 8'b1110000;
DRAM[52736] = 8'b10001100;
DRAM[52737] = 8'b10001110;
DRAM[52738] = 8'b10010000;
DRAM[52739] = 8'b10010010;
DRAM[52740] = 8'b10010100;
DRAM[52741] = 8'b10010101;
DRAM[52742] = 8'b10010101;
DRAM[52743] = 8'b10010101;
DRAM[52744] = 8'b10010110;
DRAM[52745] = 8'b10010110;
DRAM[52746] = 8'b10010110;
DRAM[52747] = 8'b10010101;
DRAM[52748] = 8'b10010101;
DRAM[52749] = 8'b10010100;
DRAM[52750] = 8'b10010100;
DRAM[52751] = 8'b10010100;
DRAM[52752] = 8'b10010101;
DRAM[52753] = 8'b10010101;
DRAM[52754] = 8'b10010110;
DRAM[52755] = 8'b10010110;
DRAM[52756] = 8'b10011000;
DRAM[52757] = 8'b10011100;
DRAM[52758] = 8'b10100010;
DRAM[52759] = 8'b10100111;
DRAM[52760] = 8'b10111111;
DRAM[52761] = 8'b11011110;
DRAM[52762] = 8'b11111010;
DRAM[52763] = 8'b11111111;
DRAM[52764] = 8'b11111100;
DRAM[52765] = 8'b11111101;
DRAM[52766] = 8'b11111111;
DRAM[52767] = 8'b11111110;
DRAM[52768] = 8'b11111110;
DRAM[52769] = 8'b11111101;
DRAM[52770] = 8'b11111010;
DRAM[52771] = 8'b11110111;
DRAM[52772] = 8'b11110101;
DRAM[52773] = 8'b11110011;
DRAM[52774] = 8'b11110011;
DRAM[52775] = 8'b11110011;
DRAM[52776] = 8'b11110010;
DRAM[52777] = 8'b11110001;
DRAM[52778] = 8'b11110001;
DRAM[52779] = 8'b11110001;
DRAM[52780] = 8'b11110010;
DRAM[52781] = 8'b11110000;
DRAM[52782] = 8'b11101101;
DRAM[52783] = 8'b11101010;
DRAM[52784] = 8'b11101100;
DRAM[52785] = 8'b11101001;
DRAM[52786] = 8'b11100110;
DRAM[52787] = 8'b11100010;
DRAM[52788] = 8'b11011110;
DRAM[52789] = 8'b11011000;
DRAM[52790] = 8'b11010000;
DRAM[52791] = 8'b11001011;
DRAM[52792] = 8'b11001110;
DRAM[52793] = 8'b11001001;
DRAM[52794] = 8'b11000110;
DRAM[52795] = 8'b11001000;
DRAM[52796] = 8'b11000111;
DRAM[52797] = 8'b11000000;
DRAM[52798] = 8'b10111100;
DRAM[52799] = 8'b10111110;
DRAM[52800] = 8'b11001000;
DRAM[52801] = 8'b11000011;
DRAM[52802] = 8'b11000000;
DRAM[52803] = 8'b10111111;
DRAM[52804] = 8'b10111101;
DRAM[52805] = 8'b10111001;
DRAM[52806] = 8'b10111001;
DRAM[52807] = 8'b10111101;
DRAM[52808] = 8'b10110000;
DRAM[52809] = 8'b10101010;
DRAM[52810] = 8'b10100011;
DRAM[52811] = 8'b10100011;
DRAM[52812] = 8'b10101010;
DRAM[52813] = 8'b10101111;
DRAM[52814] = 8'b10100111;
DRAM[52815] = 8'b10011011;
DRAM[52816] = 8'b10011100;
DRAM[52817] = 8'b10011001;
DRAM[52818] = 8'b10010110;
DRAM[52819] = 8'b10010100;
DRAM[52820] = 8'b10010100;
DRAM[52821] = 8'b10010100;
DRAM[52822] = 8'b10010011;
DRAM[52823] = 8'b10010001;
DRAM[52824] = 8'b10001110;
DRAM[52825] = 8'b10010011;
DRAM[52826] = 8'b10100000;
DRAM[52827] = 8'b10001001;
DRAM[52828] = 8'b10010000;
DRAM[52829] = 8'b10000100;
DRAM[52830] = 8'b10001110;
DRAM[52831] = 8'b10000011;
DRAM[52832] = 8'b1111011;
DRAM[52833] = 8'b1101010;
DRAM[52834] = 8'b1011101;
DRAM[52835] = 8'b1010110;
DRAM[52836] = 8'b1011001;
DRAM[52837] = 8'b1101101;
DRAM[52838] = 8'b1111011;
DRAM[52839] = 8'b1110110;
DRAM[52840] = 8'b1110011;
DRAM[52841] = 8'b1110100;
DRAM[52842] = 8'b1110010;
DRAM[52843] = 8'b1101110;
DRAM[52844] = 8'b1101100;
DRAM[52845] = 8'b1101011;
DRAM[52846] = 8'b1100101;
DRAM[52847] = 8'b1011101;
DRAM[52848] = 8'b1100111;
DRAM[52849] = 8'b1101010;
DRAM[52850] = 8'b1100011;
DRAM[52851] = 8'b1011111;
DRAM[52852] = 8'b1100110;
DRAM[52853] = 8'b1100101;
DRAM[52854] = 8'b1100000;
DRAM[52855] = 8'b1100010;
DRAM[52856] = 8'b1100110;
DRAM[52857] = 8'b1100100;
DRAM[52858] = 8'b1100100;
DRAM[52859] = 8'b1100100;
DRAM[52860] = 8'b1100011;
DRAM[52861] = 8'b1011110;
DRAM[52862] = 8'b1010100;
DRAM[52863] = 8'b1001100;
DRAM[52864] = 8'b1011011;
DRAM[52865] = 8'b1100000;
DRAM[52866] = 8'b1010011;
DRAM[52867] = 8'b1010100;
DRAM[52868] = 8'b1010100;
DRAM[52869] = 8'b1010100;
DRAM[52870] = 8'b1100001;
DRAM[52871] = 8'b1011100;
DRAM[52872] = 8'b1100000;
DRAM[52873] = 8'b1011101;
DRAM[52874] = 8'b1011110;
DRAM[52875] = 8'b1100001;
DRAM[52876] = 8'b1100010;
DRAM[52877] = 8'b1011111;
DRAM[52878] = 8'b1011111;
DRAM[52879] = 8'b1100010;
DRAM[52880] = 8'b1100110;
DRAM[52881] = 8'b1011110;
DRAM[52882] = 8'b1100000;
DRAM[52883] = 8'b1101110;
DRAM[52884] = 8'b1110010;
DRAM[52885] = 8'b1101011;
DRAM[52886] = 8'b1101100;
DRAM[52887] = 8'b1110101;
DRAM[52888] = 8'b1110110;
DRAM[52889] = 8'b1101101;
DRAM[52890] = 8'b1101101;
DRAM[52891] = 8'b1111010;
DRAM[52892] = 8'b1111110;
DRAM[52893] = 8'b1110111;
DRAM[52894] = 8'b1111000;
DRAM[52895] = 8'b10000010;
DRAM[52896] = 8'b1111110;
DRAM[52897] = 8'b10000100;
DRAM[52898] = 8'b10001010;
DRAM[52899] = 8'b10001101;
DRAM[52900] = 8'b10010001;
DRAM[52901] = 8'b10010111;
DRAM[52902] = 8'b10011111;
DRAM[52903] = 8'b10100011;
DRAM[52904] = 8'b10100011;
DRAM[52905] = 8'b10101000;
DRAM[52906] = 8'b10101101;
DRAM[52907] = 8'b10101101;
DRAM[52908] = 8'b10101011;
DRAM[52909] = 8'b10101000;
DRAM[52910] = 8'b10101001;
DRAM[52911] = 8'b10101010;
DRAM[52912] = 8'b10101110;
DRAM[52913] = 8'b10110000;
DRAM[52914] = 8'b10111001;
DRAM[52915] = 8'b11000101;
DRAM[52916] = 8'b11001101;
DRAM[52917] = 8'b11010001;
DRAM[52918] = 8'b11011001;
DRAM[52919] = 8'b11100001;
DRAM[52920] = 8'b11100010;
DRAM[52921] = 8'b11011010;
DRAM[52922] = 8'b11010010;
DRAM[52923] = 8'b11010011;
DRAM[52924] = 8'b11011011;
DRAM[52925] = 8'b11100110;
DRAM[52926] = 8'b11101100;
DRAM[52927] = 8'b11101111;
DRAM[52928] = 8'b11100101;
DRAM[52929] = 8'b11100001;
DRAM[52930] = 8'b11010111;
DRAM[52931] = 8'b11000111;
DRAM[52932] = 8'b10110101;
DRAM[52933] = 8'b10101100;
DRAM[52934] = 8'b10101100;
DRAM[52935] = 8'b10101111;
DRAM[52936] = 8'b10100000;
DRAM[52937] = 8'b10010011;
DRAM[52938] = 8'b10000110;
DRAM[52939] = 8'b10000000;
DRAM[52940] = 8'b1111101;
DRAM[52941] = 8'b1111011;
DRAM[52942] = 8'b1111011;
DRAM[52943] = 8'b1111110;
DRAM[52944] = 8'b1111001;
DRAM[52945] = 8'b1110111;
DRAM[52946] = 8'b1110101;
DRAM[52947] = 8'b1110100;
DRAM[52948] = 8'b1110100;
DRAM[52949] = 8'b1110101;
DRAM[52950] = 8'b1110011;
DRAM[52951] = 8'b1110010;
DRAM[52952] = 8'b1110010;
DRAM[52953] = 8'b1101111;
DRAM[52954] = 8'b1101101;
DRAM[52955] = 8'b1101101;
DRAM[52956] = 8'b1110000;
DRAM[52957] = 8'b1110010;
DRAM[52958] = 8'b1110011;
DRAM[52959] = 8'b1110100;
DRAM[52960] = 8'b1110100;
DRAM[52961] = 8'b1110100;
DRAM[52962] = 8'b1110100;
DRAM[52963] = 8'b1110101;
DRAM[52964] = 8'b1110101;
DRAM[52965] = 8'b1110110;
DRAM[52966] = 8'b1110110;
DRAM[52967] = 8'b1110110;
DRAM[52968] = 8'b1111000;
DRAM[52969] = 8'b1110111;
DRAM[52970] = 8'b1110111;
DRAM[52971] = 8'b1110110;
DRAM[52972] = 8'b1110101;
DRAM[52973] = 8'b1110100;
DRAM[52974] = 8'b1110011;
DRAM[52975] = 8'b1110011;
DRAM[52976] = 8'b1110011;
DRAM[52977] = 8'b1110010;
DRAM[52978] = 8'b1110010;
DRAM[52979] = 8'b1110001;
DRAM[52980] = 8'b1110000;
DRAM[52981] = 8'b1101111;
DRAM[52982] = 8'b1101111;
DRAM[52983] = 8'b1101111;
DRAM[52984] = 8'b1101101;
DRAM[52985] = 8'b1101110;
DRAM[52986] = 8'b1101111;
DRAM[52987] = 8'b1110000;
DRAM[52988] = 8'b1110001;
DRAM[52989] = 8'b1110000;
DRAM[52990] = 8'b1110000;
DRAM[52991] = 8'b1101111;
DRAM[52992] = 8'b10001100;
DRAM[52993] = 8'b10001110;
DRAM[52994] = 8'b10010000;
DRAM[52995] = 8'b10010011;
DRAM[52996] = 8'b10010101;
DRAM[52997] = 8'b10010101;
DRAM[52998] = 8'b10010101;
DRAM[52999] = 8'b10010101;
DRAM[53000] = 8'b10010110;
DRAM[53001] = 8'b10010110;
DRAM[53002] = 8'b10010110;
DRAM[53003] = 8'b10010101;
DRAM[53004] = 8'b10010101;
DRAM[53005] = 8'b10010100;
DRAM[53006] = 8'b10010100;
DRAM[53007] = 8'b10010100;
DRAM[53008] = 8'b10010100;
DRAM[53009] = 8'b10010101;
DRAM[53010] = 8'b10010110;
DRAM[53011] = 8'b10011000;
DRAM[53012] = 8'b10011010;
DRAM[53013] = 8'b10011111;
DRAM[53014] = 8'b10100110;
DRAM[53015] = 8'b10101011;
DRAM[53016] = 8'b10111110;
DRAM[53017] = 8'b11011110;
DRAM[53018] = 8'b11111011;
DRAM[53019] = 8'b11111111;
DRAM[53020] = 8'b11111010;
DRAM[53021] = 8'b11111100;
DRAM[53022] = 8'b11111111;
DRAM[53023] = 8'b11111111;
DRAM[53024] = 8'b11111111;
DRAM[53025] = 8'b11111101;
DRAM[53026] = 8'b11111001;
DRAM[53027] = 8'b11110101;
DRAM[53028] = 8'b11110001;
DRAM[53029] = 8'b11101111;
DRAM[53030] = 8'b11101101;
DRAM[53031] = 8'b11101101;
DRAM[53032] = 8'b11101110;
DRAM[53033] = 8'b11101101;
DRAM[53034] = 8'b11101101;
DRAM[53035] = 8'b11101110;
DRAM[53036] = 8'b11101111;
DRAM[53037] = 8'b11101110;
DRAM[53038] = 8'b11101011;
DRAM[53039] = 8'b11101000;
DRAM[53040] = 8'b11100100;
DRAM[53041] = 8'b11100011;
DRAM[53042] = 8'b11100001;
DRAM[53043] = 8'b11011111;
DRAM[53044] = 8'b11011101;
DRAM[53045] = 8'b11011001;
DRAM[53046] = 8'b11010011;
DRAM[53047] = 8'b11001111;
DRAM[53048] = 8'b11010011;
DRAM[53049] = 8'b11001111;
DRAM[53050] = 8'b11001100;
DRAM[53051] = 8'b11001000;
DRAM[53052] = 8'b10111110;
DRAM[53053] = 8'b10110110;
DRAM[53054] = 8'b10111001;
DRAM[53055] = 8'b11000011;
DRAM[53056] = 8'b10111000;
DRAM[53057] = 8'b10111001;
DRAM[53058] = 8'b11000000;
DRAM[53059] = 8'b11001010;
DRAM[53060] = 8'b11001010;
DRAM[53061] = 8'b11000000;
DRAM[53062] = 8'b10110100;
DRAM[53063] = 8'b10101110;
DRAM[53064] = 8'b10101011;
DRAM[53065] = 8'b10110101;
DRAM[53066] = 8'b10110100;
DRAM[53067] = 8'b10100100;
DRAM[53068] = 8'b10010111;
DRAM[53069] = 8'b10010110;
DRAM[53070] = 8'b10010111;
DRAM[53071] = 8'b10010101;
DRAM[53072] = 8'b10100001;
DRAM[53073] = 8'b10100000;
DRAM[53074] = 8'b10100000;
DRAM[53075] = 8'b10100000;
DRAM[53076] = 8'b10011110;
DRAM[53077] = 8'b10011010;
DRAM[53078] = 8'b10010101;
DRAM[53079] = 8'b10010000;
DRAM[53080] = 8'b10010010;
DRAM[53081] = 8'b10010111;
DRAM[53082] = 8'b10010100;
DRAM[53083] = 8'b10001000;
DRAM[53084] = 8'b10000100;
DRAM[53085] = 8'b10000111;
DRAM[53086] = 8'b10000100;
DRAM[53087] = 8'b1111010;
DRAM[53088] = 8'b1110101;
DRAM[53089] = 8'b1101000;
DRAM[53090] = 8'b1011110;
DRAM[53091] = 8'b1011000;
DRAM[53092] = 8'b1011011;
DRAM[53093] = 8'b1101110;
DRAM[53094] = 8'b1111100;
DRAM[53095] = 8'b1110110;
DRAM[53096] = 8'b1110100;
DRAM[53097] = 8'b1111010;
DRAM[53098] = 8'b1111000;
DRAM[53099] = 8'b1101110;
DRAM[53100] = 8'b1101000;
DRAM[53101] = 8'b1101000;
DRAM[53102] = 8'b1100011;
DRAM[53103] = 8'b1011000;
DRAM[53104] = 8'b1101011;
DRAM[53105] = 8'b1101011;
DRAM[53106] = 8'b1100100;
DRAM[53107] = 8'b1100011;
DRAM[53108] = 8'b1101010;
DRAM[53109] = 8'b1100110;
DRAM[53110] = 8'b1100000;
DRAM[53111] = 8'b1100101;
DRAM[53112] = 8'b1100100;
DRAM[53113] = 8'b1100011;
DRAM[53114] = 8'b1100010;
DRAM[53115] = 8'b1100011;
DRAM[53116] = 8'b1100011;
DRAM[53117] = 8'b1011110;
DRAM[53118] = 8'b1010101;
DRAM[53119] = 8'b1001110;
DRAM[53120] = 8'b1011010;
DRAM[53121] = 8'b1011111;
DRAM[53122] = 8'b1010100;
DRAM[53123] = 8'b1010111;
DRAM[53124] = 8'b1011001;
DRAM[53125] = 8'b1011001;
DRAM[53126] = 8'b1101000;
DRAM[53127] = 8'b1100101;
DRAM[53128] = 8'b1010111;
DRAM[53129] = 8'b1010111;
DRAM[53130] = 8'b1011011;
DRAM[53131] = 8'b1100001;
DRAM[53132] = 8'b1100001;
DRAM[53133] = 8'b1011101;
DRAM[53134] = 8'b1011101;
DRAM[53135] = 8'b1100000;
DRAM[53136] = 8'b1100111;
DRAM[53137] = 8'b1100010;
DRAM[53138] = 8'b1100001;
DRAM[53139] = 8'b1100111;
DRAM[53140] = 8'b1101111;
DRAM[53141] = 8'b1110011;
DRAM[53142] = 8'b1110010;
DRAM[53143] = 8'b1110001;
DRAM[53144] = 8'b10000001;
DRAM[53145] = 8'b1110001;
DRAM[53146] = 8'b1110001;
DRAM[53147] = 8'b10000011;
DRAM[53148] = 8'b10000111;
DRAM[53149] = 8'b1111001;
DRAM[53150] = 8'b1110110;
DRAM[53151] = 8'b10000000;
DRAM[53152] = 8'b1111011;
DRAM[53153] = 8'b1111010;
DRAM[53154] = 8'b1111110;
DRAM[53155] = 8'b10000110;
DRAM[53156] = 8'b10001110;
DRAM[53157] = 8'b10010011;
DRAM[53158] = 8'b10011000;
DRAM[53159] = 8'b10011100;
DRAM[53160] = 8'b10011110;
DRAM[53161] = 8'b10100100;
DRAM[53162] = 8'b10101100;
DRAM[53163] = 8'b10110000;
DRAM[53164] = 8'b10110001;
DRAM[53165] = 8'b10101111;
DRAM[53166] = 8'b10101111;
DRAM[53167] = 8'b10101111;
DRAM[53168] = 8'b10110011;
DRAM[53169] = 8'b10110100;
DRAM[53170] = 8'b10111100;
DRAM[53171] = 8'b11000110;
DRAM[53172] = 8'b11001110;
DRAM[53173] = 8'b11010010;
DRAM[53174] = 8'b11011010;
DRAM[53175] = 8'b11100010;
DRAM[53176] = 8'b11101011;
DRAM[53177] = 8'b11100011;
DRAM[53178] = 8'b11011100;
DRAM[53179] = 8'b11011110;
DRAM[53180] = 8'b11100110;
DRAM[53181] = 8'b11101110;
DRAM[53182] = 8'b11110001;
DRAM[53183] = 8'b11110000;
DRAM[53184] = 8'b11101111;
DRAM[53185] = 8'b11101110;
DRAM[53186] = 8'b11100101;
DRAM[53187] = 8'b11010001;
DRAM[53188] = 8'b10111010;
DRAM[53189] = 8'b10101011;
DRAM[53190] = 8'b10101000;
DRAM[53191] = 8'b10101011;
DRAM[53192] = 8'b10011111;
DRAM[53193] = 8'b10010011;
DRAM[53194] = 8'b10000111;
DRAM[53195] = 8'b10000010;
DRAM[53196] = 8'b1111111;
DRAM[53197] = 8'b1111100;
DRAM[53198] = 8'b1111100;
DRAM[53199] = 8'b1111110;
DRAM[53200] = 8'b1111101;
DRAM[53201] = 8'b1111010;
DRAM[53202] = 8'b1110111;
DRAM[53203] = 8'b1110110;
DRAM[53204] = 8'b1110101;
DRAM[53205] = 8'b1110101;
DRAM[53206] = 8'b1110011;
DRAM[53207] = 8'b1110001;
DRAM[53208] = 8'b1110011;
DRAM[53209] = 8'b1110000;
DRAM[53210] = 8'b1101110;
DRAM[53211] = 8'b1101110;
DRAM[53212] = 8'b1110000;
DRAM[53213] = 8'b1110011;
DRAM[53214] = 8'b1110100;
DRAM[53215] = 8'b1110100;
DRAM[53216] = 8'b1110101;
DRAM[53217] = 8'b1110101;
DRAM[53218] = 8'b1110101;
DRAM[53219] = 8'b1110101;
DRAM[53220] = 8'b1110101;
DRAM[53221] = 8'b1110101;
DRAM[53222] = 8'b1110101;
DRAM[53223] = 8'b1110101;
DRAM[53224] = 8'b1110111;
DRAM[53225] = 8'b1110111;
DRAM[53226] = 8'b1110110;
DRAM[53227] = 8'b1110101;
DRAM[53228] = 8'b1110100;
DRAM[53229] = 8'b1110100;
DRAM[53230] = 8'b1110011;
DRAM[53231] = 8'b1110010;
DRAM[53232] = 8'b1110001;
DRAM[53233] = 8'b1110001;
DRAM[53234] = 8'b1110000;
DRAM[53235] = 8'b1101111;
DRAM[53236] = 8'b1101110;
DRAM[53237] = 8'b1101110;
DRAM[53238] = 8'b1101101;
DRAM[53239] = 8'b1101101;
DRAM[53240] = 8'b1101100;
DRAM[53241] = 8'b1101101;
DRAM[53242] = 8'b1101111;
DRAM[53243] = 8'b1110000;
DRAM[53244] = 8'b1110001;
DRAM[53245] = 8'b1110000;
DRAM[53246] = 8'b1101111;
DRAM[53247] = 8'b1101110;
DRAM[53248] = 8'b10010010;
DRAM[53249] = 8'b10010011;
DRAM[53250] = 8'b10010011;
DRAM[53251] = 8'b10010100;
DRAM[53252] = 8'b10010101;
DRAM[53253] = 8'b10010110;
DRAM[53254] = 8'b10010111;
DRAM[53255] = 8'b10011000;
DRAM[53256] = 8'b10010110;
DRAM[53257] = 8'b10010111;
DRAM[53258] = 8'b10010111;
DRAM[53259] = 8'b10010110;
DRAM[53260] = 8'b10010011;
DRAM[53261] = 8'b10010010;
DRAM[53262] = 8'b10010011;
DRAM[53263] = 8'b10010100;
DRAM[53264] = 8'b10011001;
DRAM[53265] = 8'b10010001;
DRAM[53266] = 8'b10010010;
DRAM[53267] = 8'b10011011;
DRAM[53268] = 8'b10011111;
DRAM[53269] = 8'b10011100;
DRAM[53270] = 8'b10011111;
DRAM[53271] = 8'b10101001;
DRAM[53272] = 8'b11000101;
DRAM[53273] = 8'b11100101;
DRAM[53274] = 8'b11111111;
DRAM[53275] = 8'b11111111;
DRAM[53276] = 8'b11111001;
DRAM[53277] = 8'b11111010;
DRAM[53278] = 8'b11111111;
DRAM[53279] = 8'b11111111;
DRAM[53280] = 8'b11111111;
DRAM[53281] = 8'b11111100;
DRAM[53282] = 8'b11110111;
DRAM[53283] = 8'b11110101;
DRAM[53284] = 8'b11110100;
DRAM[53285] = 8'b11110011;
DRAM[53286] = 8'b11110001;
DRAM[53287] = 8'b11110000;
DRAM[53288] = 8'b11110001;
DRAM[53289] = 8'b11110010;
DRAM[53290] = 8'b11110010;
DRAM[53291] = 8'b11110010;
DRAM[53292] = 8'b11101111;
DRAM[53293] = 8'b11101011;
DRAM[53294] = 8'b11100111;
DRAM[53295] = 8'b11100100;
DRAM[53296] = 8'b11100101;
DRAM[53297] = 8'b11100101;
DRAM[53298] = 8'b11100011;
DRAM[53299] = 8'b11100010;
DRAM[53300] = 8'b11100000;
DRAM[53301] = 8'b11011111;
DRAM[53302] = 8'b11011101;
DRAM[53303] = 8'b11011101;
DRAM[53304] = 8'b11001101;
DRAM[53305] = 8'b11000110;
DRAM[53306] = 8'b11001001;
DRAM[53307] = 8'b11010110;
DRAM[53308] = 8'b11011001;
DRAM[53309] = 8'b11001110;
DRAM[53310] = 8'b11000110;
DRAM[53311] = 8'b11000111;
DRAM[53312] = 8'b10111000;
DRAM[53313] = 8'b11000001;
DRAM[53314] = 8'b11000001;
DRAM[53315] = 8'b10110110;
DRAM[53316] = 8'b10110000;
DRAM[53317] = 8'b10110111;
DRAM[53318] = 8'b10111100;
DRAM[53319] = 8'b10111010;
DRAM[53320] = 8'b10100100;
DRAM[53321] = 8'b10100000;
DRAM[53322] = 8'b10100000;
DRAM[53323] = 8'b10100011;
DRAM[53324] = 8'b10011111;
DRAM[53325] = 8'b10010110;
DRAM[53326] = 8'b10010111;
DRAM[53327] = 8'b10100000;
DRAM[53328] = 8'b10100100;
DRAM[53329] = 8'b10011010;
DRAM[53330] = 8'b10011010;
DRAM[53331] = 8'b10011001;
DRAM[53332] = 8'b10001110;
DRAM[53333] = 8'b10001100;
DRAM[53334] = 8'b10010010;
DRAM[53335] = 8'b10010011;
DRAM[53336] = 8'b10011000;
DRAM[53337] = 8'b10010111;
DRAM[53338] = 8'b10001101;
DRAM[53339] = 8'b10001000;
DRAM[53340] = 8'b10001101;
DRAM[53341] = 8'b10001000;
DRAM[53342] = 8'b1111101;
DRAM[53343] = 8'b1111100;
DRAM[53344] = 8'b1110011;
DRAM[53345] = 8'b1011111;
DRAM[53346] = 8'b1011110;
DRAM[53347] = 8'b1011110;
DRAM[53348] = 8'b1101010;
DRAM[53349] = 8'b1110101;
DRAM[53350] = 8'b1101101;
DRAM[53351] = 8'b1110011;
DRAM[53352] = 8'b1110001;
DRAM[53353] = 8'b1101100;
DRAM[53354] = 8'b1110110;
DRAM[53355] = 8'b1101110;
DRAM[53356] = 8'b1011011;
DRAM[53357] = 8'b1101010;
DRAM[53358] = 8'b1110011;
DRAM[53359] = 8'b1010110;
DRAM[53360] = 8'b1110111;
DRAM[53361] = 8'b1101011;
DRAM[53362] = 8'b1010111;
DRAM[53363] = 8'b1011101;
DRAM[53364] = 8'b1111010;
DRAM[53365] = 8'b1011101;
DRAM[53366] = 8'b1101010;
DRAM[53367] = 8'b1100010;
DRAM[53368] = 8'b1100011;
DRAM[53369] = 8'b1101011;
DRAM[53370] = 8'b1101101;
DRAM[53371] = 8'b1100100;
DRAM[53372] = 8'b1011100;
DRAM[53373] = 8'b1011000;
DRAM[53374] = 8'b1010011;
DRAM[53375] = 8'b1001101;
DRAM[53376] = 8'b1011001;
DRAM[53377] = 8'b1011001;
DRAM[53378] = 8'b1011111;
DRAM[53379] = 8'b1011101;
DRAM[53380] = 8'b1010101;
DRAM[53381] = 8'b1011100;
DRAM[53382] = 8'b1101000;
DRAM[53383] = 8'b1100110;
DRAM[53384] = 8'b1100101;
DRAM[53385] = 8'b1010111;
DRAM[53386] = 8'b1011100;
DRAM[53387] = 8'b1101000;
DRAM[53388] = 8'b1100101;
DRAM[53389] = 8'b1100000;
DRAM[53390] = 8'b1100001;
DRAM[53391] = 8'b1100000;
DRAM[53392] = 8'b1100111;
DRAM[53393] = 8'b1100110;
DRAM[53394] = 8'b1100101;
DRAM[53395] = 8'b1100110;
DRAM[53396] = 8'b1110000;
DRAM[53397] = 8'b1111000;
DRAM[53398] = 8'b1110001;
DRAM[53399] = 8'b1100101;
DRAM[53400] = 8'b1111101;
DRAM[53401] = 8'b1110111;
DRAM[53402] = 8'b1111001;
DRAM[53403] = 8'b1101000;
DRAM[53404] = 8'b1111111;
DRAM[53405] = 8'b10000100;
DRAM[53406] = 8'b10001101;
DRAM[53407] = 8'b1111101;
DRAM[53408] = 8'b10001001;
DRAM[53409] = 8'b10001011;
DRAM[53410] = 8'b10001101;
DRAM[53411] = 8'b10001110;
DRAM[53412] = 8'b10001111;
DRAM[53413] = 8'b10010010;
DRAM[53414] = 8'b10010110;
DRAM[53415] = 8'b10011010;
DRAM[53416] = 8'b10101000;
DRAM[53417] = 8'b10101110;
DRAM[53418] = 8'b10101011;
DRAM[53419] = 8'b10101011;
DRAM[53420] = 8'b10110011;
DRAM[53421] = 8'b10110010;
DRAM[53422] = 8'b10101111;
DRAM[53423] = 8'b10110101;
DRAM[53424] = 8'b10111011;
DRAM[53425] = 8'b11000000;
DRAM[53426] = 8'b11000110;
DRAM[53427] = 8'b11001011;
DRAM[53428] = 8'b11001101;
DRAM[53429] = 8'b11010010;
DRAM[53430] = 8'b11011000;
DRAM[53431] = 8'b11011101;
DRAM[53432] = 8'b11011100;
DRAM[53433] = 8'b11100000;
DRAM[53434] = 8'b11100110;
DRAM[53435] = 8'b11101010;
DRAM[53436] = 8'b11101100;
DRAM[53437] = 8'b11101101;
DRAM[53438] = 8'b11101110;
DRAM[53439] = 8'b11101110;
DRAM[53440] = 8'b11101110;
DRAM[53441] = 8'b11101011;
DRAM[53442] = 8'b11011111;
DRAM[53443] = 8'b11001111;
DRAM[53444] = 8'b11000110;
DRAM[53445] = 8'b11000100;
DRAM[53446] = 8'b10111111;
DRAM[53447] = 8'b10111000;
DRAM[53448] = 8'b10100110;
DRAM[53449] = 8'b10011001;
DRAM[53450] = 8'b10001001;
DRAM[53451] = 8'b10000000;
DRAM[53452] = 8'b1111101;
DRAM[53453] = 8'b1111101;
DRAM[53454] = 8'b1111100;
DRAM[53455] = 8'b1111001;
DRAM[53456] = 8'b1110110;
DRAM[53457] = 8'b1111001;
DRAM[53458] = 8'b1111000;
DRAM[53459] = 8'b1110100;
DRAM[53460] = 8'b1110011;
DRAM[53461] = 8'b1110110;
DRAM[53462] = 8'b1110111;
DRAM[53463] = 8'b1110100;
DRAM[53464] = 8'b1110010;
DRAM[53465] = 8'b1110001;
DRAM[53466] = 8'b1110000;
DRAM[53467] = 8'b1101110;
DRAM[53468] = 8'b1101110;
DRAM[53469] = 8'b1101111;
DRAM[53470] = 8'b1110000;
DRAM[53471] = 8'b1110001;
DRAM[53472] = 8'b1110101;
DRAM[53473] = 8'b1110101;
DRAM[53474] = 8'b1110100;
DRAM[53475] = 8'b1110011;
DRAM[53476] = 8'b1110011;
DRAM[53477] = 8'b1110100;
DRAM[53478] = 8'b1110100;
DRAM[53479] = 8'b1110101;
DRAM[53480] = 8'b1110101;
DRAM[53481] = 8'b1110101;
DRAM[53482] = 8'b1110101;
DRAM[53483] = 8'b1110101;
DRAM[53484] = 8'b1110100;
DRAM[53485] = 8'b1110011;
DRAM[53486] = 8'b1110010;
DRAM[53487] = 8'b1110001;
DRAM[53488] = 8'b1110001;
DRAM[53489] = 8'b1110010;
DRAM[53490] = 8'b1110010;
DRAM[53491] = 8'b1110001;
DRAM[53492] = 8'b1110000;
DRAM[53493] = 8'b1101111;
DRAM[53494] = 8'b1101110;
DRAM[53495] = 8'b1101101;
DRAM[53496] = 8'b1101101;
DRAM[53497] = 8'b1101101;
DRAM[53498] = 8'b1101110;
DRAM[53499] = 8'b1101111;
DRAM[53500] = 8'b1110000;
DRAM[53501] = 8'b1110000;
DRAM[53502] = 8'b1110001;
DRAM[53503] = 8'b1110001;
DRAM[53504] = 8'b10010100;
DRAM[53505] = 8'b10010100;
DRAM[53506] = 8'b10010100;
DRAM[53507] = 8'b10010101;
DRAM[53508] = 8'b10010110;
DRAM[53509] = 8'b10010110;
DRAM[53510] = 8'b10010111;
DRAM[53511] = 8'b10010111;
DRAM[53512] = 8'b10010111;
DRAM[53513] = 8'b10011000;
DRAM[53514] = 8'b10011001;
DRAM[53515] = 8'b10010111;
DRAM[53516] = 8'b10010101;
DRAM[53517] = 8'b10010011;
DRAM[53518] = 8'b10010100;
DRAM[53519] = 8'b10010101;
DRAM[53520] = 8'b10011000;
DRAM[53521] = 8'b10010100;
DRAM[53522] = 8'b10010111;
DRAM[53523] = 8'b10100000;
DRAM[53524] = 8'b10100100;
DRAM[53525] = 8'b10100100;
DRAM[53526] = 8'b10101111;
DRAM[53527] = 8'b10111101;
DRAM[53528] = 8'b11011001;
DRAM[53529] = 8'b11101110;
DRAM[53530] = 8'b11111110;
DRAM[53531] = 8'b11111101;
DRAM[53532] = 8'b11111010;
DRAM[53533] = 8'b11111101;
DRAM[53534] = 8'b11111111;
DRAM[53535] = 8'b11111101;
DRAM[53536] = 8'b11111000;
DRAM[53537] = 8'b11110110;
DRAM[53538] = 8'b11110101;
DRAM[53539] = 8'b11110110;
DRAM[53540] = 8'b11111000;
DRAM[53541] = 8'b11111010;
DRAM[53542] = 8'b11111010;
DRAM[53543] = 8'b11111001;
DRAM[53544] = 8'b11101101;
DRAM[53545] = 8'b11101100;
DRAM[53546] = 8'b11101011;
DRAM[53547] = 8'b11101001;
DRAM[53548] = 8'b11100111;
DRAM[53549] = 8'b11100101;
DRAM[53550] = 8'b11100100;
DRAM[53551] = 8'b11100011;
DRAM[53552] = 8'b11100011;
DRAM[53553] = 8'b11100011;
DRAM[53554] = 8'b11100010;
DRAM[53555] = 8'b11100001;
DRAM[53556] = 8'b11011111;
DRAM[53557] = 8'b11011110;
DRAM[53558] = 8'b11011101;
DRAM[53559] = 8'b11011100;
DRAM[53560] = 8'b11011001;
DRAM[53561] = 8'b11010101;
DRAM[53562] = 8'b11001110;
DRAM[53563] = 8'b11001001;
DRAM[53564] = 8'b11001001;
DRAM[53565] = 8'b11001011;
DRAM[53566] = 8'b11001000;
DRAM[53567] = 8'b11000100;
DRAM[53568] = 8'b11001001;
DRAM[53569] = 8'b11001110;
DRAM[53570] = 8'b11001000;
DRAM[53571] = 8'b10110111;
DRAM[53572] = 8'b10101100;
DRAM[53573] = 8'b10101101;
DRAM[53574] = 8'b10101110;
DRAM[53575] = 8'b10101010;
DRAM[53576] = 8'b10101100;
DRAM[53577] = 8'b10101100;
DRAM[53578] = 8'b10100110;
DRAM[53579] = 8'b10011011;
DRAM[53580] = 8'b10010110;
DRAM[53581] = 8'b10011010;
DRAM[53582] = 8'b10100010;
DRAM[53583] = 8'b10100110;
DRAM[53584] = 8'b10101011;
DRAM[53585] = 8'b10011100;
DRAM[53586] = 8'b10011000;
DRAM[53587] = 8'b10011000;
DRAM[53588] = 8'b10010011;
DRAM[53589] = 8'b10010101;
DRAM[53590] = 8'b10011100;
DRAM[53591] = 8'b10011010;
DRAM[53592] = 8'b10010111;
DRAM[53593] = 8'b10010011;
DRAM[53594] = 8'b10010000;
DRAM[53595] = 8'b10001011;
DRAM[53596] = 8'b10000110;
DRAM[53597] = 8'b10000100;
DRAM[53598] = 8'b10000100;
DRAM[53599] = 8'b10000011;
DRAM[53600] = 8'b1110001;
DRAM[53601] = 8'b1100011;
DRAM[53602] = 8'b1100100;
DRAM[53603] = 8'b1011111;
DRAM[53604] = 8'b1101001;
DRAM[53605] = 8'b1111000;
DRAM[53606] = 8'b1110001;
DRAM[53607] = 8'b1110101;
DRAM[53608] = 8'b1110000;
DRAM[53609] = 8'b1101111;
DRAM[53610] = 8'b1110100;
DRAM[53611] = 8'b1101100;
DRAM[53612] = 8'b1011111;
DRAM[53613] = 8'b1101010;
DRAM[53614] = 8'b1101101;
DRAM[53615] = 8'b1010110;
DRAM[53616] = 8'b1101101;
DRAM[53617] = 8'b1101011;
DRAM[53618] = 8'b1011101;
DRAM[53619] = 8'b1011101;
DRAM[53620] = 8'b1110010;
DRAM[53621] = 8'b1011010;
DRAM[53622] = 8'b1101000;
DRAM[53623] = 8'b1100100;
DRAM[53624] = 8'b1100111;
DRAM[53625] = 8'b1101000;
DRAM[53626] = 8'b1100110;
DRAM[53627] = 8'b1100001;
DRAM[53628] = 8'b1011111;
DRAM[53629] = 8'b1011110;
DRAM[53630] = 8'b1010110;
DRAM[53631] = 8'b1001011;
DRAM[53632] = 8'b1011001;
DRAM[53633] = 8'b1011001;
DRAM[53634] = 8'b1100000;
DRAM[53635] = 8'b1011111;
DRAM[53636] = 8'b1010111;
DRAM[53637] = 8'b1011101;
DRAM[53638] = 8'b1100111;
DRAM[53639] = 8'b1100100;
DRAM[53640] = 8'b1100011;
DRAM[53641] = 8'b1100001;
DRAM[53642] = 8'b1101000;
DRAM[53643] = 8'b1101000;
DRAM[53644] = 8'b1100010;
DRAM[53645] = 8'b1100110;
DRAM[53646] = 8'b1101011;
DRAM[53647] = 8'b1100110;
DRAM[53648] = 8'b1100011;
DRAM[53649] = 8'b1101000;
DRAM[53650] = 8'b1101011;
DRAM[53651] = 8'b1101000;
DRAM[53652] = 8'b1101001;
DRAM[53653] = 8'b1101110;
DRAM[53654] = 8'b1110001;
DRAM[53655] = 8'b1101111;
DRAM[53656] = 8'b1111010;
DRAM[53657] = 8'b1111110;
DRAM[53658] = 8'b1110110;
DRAM[53659] = 8'b1110000;
DRAM[53660] = 8'b1110001;
DRAM[53661] = 8'b10000001;
DRAM[53662] = 8'b10000101;
DRAM[53663] = 8'b10000100;
DRAM[53664] = 8'b10000011;
DRAM[53665] = 8'b10000101;
DRAM[53666] = 8'b10001000;
DRAM[53667] = 8'b10001011;
DRAM[53668] = 8'b10001101;
DRAM[53669] = 8'b10010001;
DRAM[53670] = 8'b10010111;
DRAM[53671] = 8'b10011010;
DRAM[53672] = 8'b10011010;
DRAM[53673] = 8'b10100011;
DRAM[53674] = 8'b10100101;
DRAM[53675] = 8'b10101001;
DRAM[53676] = 8'b10110101;
DRAM[53677] = 8'b10110111;
DRAM[53678] = 8'b10110110;
DRAM[53679] = 8'b10111100;
DRAM[53680] = 8'b10111011;
DRAM[53681] = 8'b10111110;
DRAM[53682] = 8'b11000100;
DRAM[53683] = 8'b11001001;
DRAM[53684] = 8'b11001110;
DRAM[53685] = 8'b11010100;
DRAM[53686] = 8'b11011001;
DRAM[53687] = 8'b11011101;
DRAM[53688] = 8'b11100001;
DRAM[53689] = 8'b11100110;
DRAM[53690] = 8'b11101100;
DRAM[53691] = 8'b11101110;
DRAM[53692] = 8'b11101100;
DRAM[53693] = 8'b11101010;
DRAM[53694] = 8'b11101011;
DRAM[53695] = 8'b11101110;
DRAM[53696] = 8'b11110001;
DRAM[53697] = 8'b11100000;
DRAM[53698] = 8'b11000111;
DRAM[53699] = 8'b10111000;
DRAM[53700] = 8'b10111011;
DRAM[53701] = 8'b10111111;
DRAM[53702] = 8'b10110111;
DRAM[53703] = 8'b10101001;
DRAM[53704] = 8'b10101011;
DRAM[53705] = 8'b10100100;
DRAM[53706] = 8'b10011000;
DRAM[53707] = 8'b10001100;
DRAM[53708] = 8'b10000011;
DRAM[53709] = 8'b1111101;
DRAM[53710] = 8'b1111011;
DRAM[53711] = 8'b1111001;
DRAM[53712] = 8'b1110111;
DRAM[53713] = 8'b1111001;
DRAM[53714] = 8'b1111000;
DRAM[53715] = 8'b1110100;
DRAM[53716] = 8'b1110100;
DRAM[53717] = 8'b1110111;
DRAM[53718] = 8'b1110111;
DRAM[53719] = 8'b1110101;
DRAM[53720] = 8'b1110011;
DRAM[53721] = 8'b1110010;
DRAM[53722] = 8'b1110000;
DRAM[53723] = 8'b1101111;
DRAM[53724] = 8'b1101110;
DRAM[53725] = 8'b1101111;
DRAM[53726] = 8'b1110000;
DRAM[53727] = 8'b1110001;
DRAM[53728] = 8'b1110101;
DRAM[53729] = 8'b1110100;
DRAM[53730] = 8'b1110100;
DRAM[53731] = 8'b1110011;
DRAM[53732] = 8'b1110011;
DRAM[53733] = 8'b1110011;
DRAM[53734] = 8'b1110100;
DRAM[53735] = 8'b1110100;
DRAM[53736] = 8'b1110110;
DRAM[53737] = 8'b1110110;
DRAM[53738] = 8'b1110110;
DRAM[53739] = 8'b1110110;
DRAM[53740] = 8'b1110101;
DRAM[53741] = 8'b1110011;
DRAM[53742] = 8'b1110010;
DRAM[53743] = 8'b1110001;
DRAM[53744] = 8'b1110001;
DRAM[53745] = 8'b1110001;
DRAM[53746] = 8'b1110001;
DRAM[53747] = 8'b1110001;
DRAM[53748] = 8'b1110000;
DRAM[53749] = 8'b1101111;
DRAM[53750] = 8'b1101110;
DRAM[53751] = 8'b1101101;
DRAM[53752] = 8'b1101101;
DRAM[53753] = 8'b1101101;
DRAM[53754] = 8'b1101110;
DRAM[53755] = 8'b1101110;
DRAM[53756] = 8'b1101111;
DRAM[53757] = 8'b1110000;
DRAM[53758] = 8'b1110001;
DRAM[53759] = 8'b1110001;
DRAM[53760] = 8'b10010110;
DRAM[53761] = 8'b10010110;
DRAM[53762] = 8'b10010110;
DRAM[53763] = 8'b10010110;
DRAM[53764] = 8'b10010110;
DRAM[53765] = 8'b10010110;
DRAM[53766] = 8'b10010111;
DRAM[53767] = 8'b10010111;
DRAM[53768] = 8'b10011001;
DRAM[53769] = 8'b10011010;
DRAM[53770] = 8'b10011011;
DRAM[53771] = 8'b10011001;
DRAM[53772] = 8'b10010111;
DRAM[53773] = 8'b10010110;
DRAM[53774] = 8'b10010110;
DRAM[53775] = 8'b10010111;
DRAM[53776] = 8'b10011001;
DRAM[53777] = 8'b10011000;
DRAM[53778] = 8'b10011100;
DRAM[53779] = 8'b10100001;
DRAM[53780] = 8'b10100100;
DRAM[53781] = 8'b10101010;
DRAM[53782] = 8'b10111110;
DRAM[53783] = 8'b11010011;
DRAM[53784] = 8'b11101111;
DRAM[53785] = 8'b11111001;
DRAM[53786] = 8'b11111101;
DRAM[53787] = 8'b11111011;
DRAM[53788] = 8'b11111100;
DRAM[53789] = 8'b11111111;
DRAM[53790] = 8'b11111111;
DRAM[53791] = 8'b11111001;
DRAM[53792] = 8'b11111001;
DRAM[53793] = 8'b11111000;
DRAM[53794] = 8'b11110110;
DRAM[53795] = 8'b11110111;
DRAM[53796] = 8'b11110111;
DRAM[53797] = 8'b11110111;
DRAM[53798] = 8'b11110100;
DRAM[53799] = 8'b11110010;
DRAM[53800] = 8'b11110000;
DRAM[53801] = 8'b11101110;
DRAM[53802] = 8'b11101011;
DRAM[53803] = 8'b11101000;
DRAM[53804] = 8'b11100111;
DRAM[53805] = 8'b11100111;
DRAM[53806] = 8'b11101000;
DRAM[53807] = 8'b11101001;
DRAM[53808] = 8'b11100011;
DRAM[53809] = 8'b11100010;
DRAM[53810] = 8'b11100001;
DRAM[53811] = 8'b11011111;
DRAM[53812] = 8'b11011110;
DRAM[53813] = 8'b11011100;
DRAM[53814] = 8'b11011011;
DRAM[53815] = 8'b11011010;
DRAM[53816] = 8'b11011001;
DRAM[53817] = 8'b11011010;
DRAM[53818] = 8'b11001111;
DRAM[53819] = 8'b10111111;
DRAM[53820] = 8'b10111110;
DRAM[53821] = 8'b11001000;
DRAM[53822] = 8'b11001000;
DRAM[53823] = 8'b10111111;
DRAM[53824] = 8'b10111101;
DRAM[53825] = 8'b11000000;
DRAM[53826] = 8'b10111010;
DRAM[53827] = 8'b10101010;
DRAM[53828] = 8'b10100001;
DRAM[53829] = 8'b10100011;
DRAM[53830] = 8'b10100101;
DRAM[53831] = 8'b10100010;
DRAM[53832] = 8'b10110000;
DRAM[53833] = 8'b10110100;
DRAM[53834] = 8'b10101100;
DRAM[53835] = 8'b10011011;
DRAM[53836] = 8'b10010111;
DRAM[53837] = 8'b10100011;
DRAM[53838] = 8'b10101010;
DRAM[53839] = 8'b10100111;
DRAM[53840] = 8'b10101001;
DRAM[53841] = 8'b10011010;
DRAM[53842] = 8'b10010111;
DRAM[53843] = 8'b10011100;
DRAM[53844] = 8'b10011011;
DRAM[53845] = 8'b10011101;
DRAM[53846] = 8'b10011110;
DRAM[53847] = 8'b10011000;
DRAM[53848] = 8'b10011000;
DRAM[53849] = 8'b10001110;
DRAM[53850] = 8'b10010011;
DRAM[53851] = 8'b10010000;
DRAM[53852] = 8'b1111110;
DRAM[53853] = 8'b10000000;
DRAM[53854] = 8'b10001011;
DRAM[53855] = 8'b10000110;
DRAM[53856] = 8'b1101111;
DRAM[53857] = 8'b1101010;
DRAM[53858] = 8'b1101101;
DRAM[53859] = 8'b1100010;
DRAM[53860] = 8'b1101001;
DRAM[53861] = 8'b1111100;
DRAM[53862] = 8'b1111000;
DRAM[53863] = 8'b1111001;
DRAM[53864] = 8'b1110000;
DRAM[53865] = 8'b1110101;
DRAM[53866] = 8'b1110010;
DRAM[53867] = 8'b1101000;
DRAM[53868] = 8'b1100101;
DRAM[53869] = 8'b1101011;
DRAM[53870] = 8'b1101000;
DRAM[53871] = 8'b1011100;
DRAM[53872] = 8'b1100001;
DRAM[53873] = 8'b1101001;
DRAM[53874] = 8'b1100010;
DRAM[53875] = 8'b1011100;
DRAM[53876] = 8'b1100111;
DRAM[53877] = 8'b1011001;
DRAM[53878] = 8'b1100101;
DRAM[53879] = 8'b1100110;
DRAM[53880] = 8'b1101010;
DRAM[53881] = 8'b1100100;
DRAM[53882] = 8'b1011110;
DRAM[53883] = 8'b1011101;
DRAM[53884] = 8'b1100010;
DRAM[53885] = 8'b1100011;
DRAM[53886] = 8'b1011000;
DRAM[53887] = 8'b1001011;
DRAM[53888] = 8'b1011001;
DRAM[53889] = 8'b1011010;
DRAM[53890] = 8'b1100010;
DRAM[53891] = 8'b1100010;
DRAM[53892] = 8'b1011010;
DRAM[53893] = 8'b1100000;
DRAM[53894] = 8'b1100111;
DRAM[53895] = 8'b1100001;
DRAM[53896] = 8'b1011011;
DRAM[53897] = 8'b1100011;
DRAM[53898] = 8'b1101011;
DRAM[53899] = 8'b1100100;
DRAM[53900] = 8'b1011100;
DRAM[53901] = 8'b1100111;
DRAM[53902] = 8'b1101111;
DRAM[53903] = 8'b1100101;
DRAM[53904] = 8'b1100111;
DRAM[53905] = 8'b1101001;
DRAM[53906] = 8'b1101001;
DRAM[53907] = 8'b1100101;
DRAM[53908] = 8'b1100110;
DRAM[53909] = 8'b1101101;
DRAM[53910] = 8'b1110010;
DRAM[53911] = 8'b1110100;
DRAM[53912] = 8'b1110110;
DRAM[53913] = 8'b10000100;
DRAM[53914] = 8'b1111010;
DRAM[53915] = 8'b1111110;
DRAM[53916] = 8'b1101001;
DRAM[53917] = 8'b1111100;
DRAM[53918] = 8'b1110111;
DRAM[53919] = 8'b1111110;
DRAM[53920] = 8'b10000101;
DRAM[53921] = 8'b10001000;
DRAM[53922] = 8'b10001011;
DRAM[53923] = 8'b10001110;
DRAM[53924] = 8'b10010000;
DRAM[53925] = 8'b10010011;
DRAM[53926] = 8'b10011000;
DRAM[53927] = 8'b10011011;
DRAM[53928] = 8'b10010111;
DRAM[53929] = 8'b10100001;
DRAM[53930] = 8'b10100100;
DRAM[53931] = 8'b10101001;
DRAM[53932] = 8'b10110101;
DRAM[53933] = 8'b10110111;
DRAM[53934] = 8'b10110100;
DRAM[53935] = 8'b10111010;
DRAM[53936] = 8'b10111010;
DRAM[53937] = 8'b10111011;
DRAM[53938] = 8'b10111111;
DRAM[53939] = 8'b11000101;
DRAM[53940] = 8'b11001101;
DRAM[53941] = 8'b11010011;
DRAM[53942] = 8'b11010111;
DRAM[53943] = 8'b11011000;
DRAM[53944] = 8'b11011111;
DRAM[53945] = 8'b11100101;
DRAM[53946] = 8'b11101011;
DRAM[53947] = 8'b11101100;
DRAM[53948] = 8'b11101001;
DRAM[53949] = 8'b11101000;
DRAM[53950] = 8'b11101011;
DRAM[53951] = 8'b11101111;
DRAM[53952] = 8'b11110010;
DRAM[53953] = 8'b11101001;
DRAM[53954] = 8'b11010111;
DRAM[53955] = 8'b11000010;
DRAM[53956] = 8'b10110011;
DRAM[53957] = 8'b10101001;
DRAM[53958] = 8'b10011111;
DRAM[53959] = 8'b10011000;
DRAM[53960] = 8'b10010110;
DRAM[53961] = 8'b10010101;
DRAM[53962] = 8'b10010001;
DRAM[53963] = 8'b10001001;
DRAM[53964] = 8'b10000001;
DRAM[53965] = 8'b1111101;
DRAM[53966] = 8'b1111101;
DRAM[53967] = 8'b1111111;
DRAM[53968] = 8'b1110111;
DRAM[53969] = 8'b1111010;
DRAM[53970] = 8'b1111001;
DRAM[53971] = 8'b1110101;
DRAM[53972] = 8'b1110100;
DRAM[53973] = 8'b1110111;
DRAM[53974] = 8'b1111000;
DRAM[53975] = 8'b1110101;
DRAM[53976] = 8'b1110011;
DRAM[53977] = 8'b1110010;
DRAM[53978] = 8'b1110000;
DRAM[53979] = 8'b1101111;
DRAM[53980] = 8'b1101111;
DRAM[53981] = 8'b1101111;
DRAM[53982] = 8'b1110000;
DRAM[53983] = 8'b1110001;
DRAM[53984] = 8'b1110100;
DRAM[53985] = 8'b1110011;
DRAM[53986] = 8'b1110011;
DRAM[53987] = 8'b1110010;
DRAM[53988] = 8'b1110010;
DRAM[53989] = 8'b1110011;
DRAM[53990] = 8'b1110100;
DRAM[53991] = 8'b1110100;
DRAM[53992] = 8'b1110110;
DRAM[53993] = 8'b1110110;
DRAM[53994] = 8'b1110110;
DRAM[53995] = 8'b1110110;
DRAM[53996] = 8'b1110101;
DRAM[53997] = 8'b1110100;
DRAM[53998] = 8'b1110011;
DRAM[53999] = 8'b1110010;
DRAM[54000] = 8'b1110000;
DRAM[54001] = 8'b1110001;
DRAM[54002] = 8'b1110001;
DRAM[54003] = 8'b1110000;
DRAM[54004] = 8'b1110000;
DRAM[54005] = 8'b1101110;
DRAM[54006] = 8'b1101101;
DRAM[54007] = 8'b1101100;
DRAM[54008] = 8'b1101100;
DRAM[54009] = 8'b1101100;
DRAM[54010] = 8'b1101101;
DRAM[54011] = 8'b1101110;
DRAM[54012] = 8'b1101111;
DRAM[54013] = 8'b1101111;
DRAM[54014] = 8'b1110000;
DRAM[54015] = 8'b1110000;
DRAM[54016] = 8'b10011000;
DRAM[54017] = 8'b10011000;
DRAM[54018] = 8'b10011000;
DRAM[54019] = 8'b10010111;
DRAM[54020] = 8'b10010111;
DRAM[54021] = 8'b10010111;
DRAM[54022] = 8'b10010111;
DRAM[54023] = 8'b10010111;
DRAM[54024] = 8'b10011011;
DRAM[54025] = 8'b10011100;
DRAM[54026] = 8'b10011101;
DRAM[54027] = 8'b10011100;
DRAM[54028] = 8'b10011001;
DRAM[54029] = 8'b10011000;
DRAM[54030] = 8'b10011000;
DRAM[54031] = 8'b10011001;
DRAM[54032] = 8'b10011010;
DRAM[54033] = 8'b10011010;
DRAM[54034] = 8'b10011011;
DRAM[54035] = 8'b10011100;
DRAM[54036] = 8'b10011110;
DRAM[54037] = 8'b10101010;
DRAM[54038] = 8'b11000111;
DRAM[54039] = 8'b11100010;
DRAM[54040] = 8'b11111010;
DRAM[54041] = 8'b11111110;
DRAM[54042] = 8'b11111111;
DRAM[54043] = 8'b11111100;
DRAM[54044] = 8'b11111101;
DRAM[54045] = 8'b11111111;
DRAM[54046] = 8'b11111101;
DRAM[54047] = 8'b11110110;
DRAM[54048] = 8'b11111110;
DRAM[54049] = 8'b11111100;
DRAM[54050] = 8'b11111011;
DRAM[54051] = 8'b11111010;
DRAM[54052] = 8'b11111000;
DRAM[54053] = 8'b11110101;
DRAM[54054] = 8'b11110001;
DRAM[54055] = 8'b11101101;
DRAM[54056] = 8'b11101111;
DRAM[54057] = 8'b11101101;
DRAM[54058] = 8'b11101011;
DRAM[54059] = 8'b11101010;
DRAM[54060] = 8'b11101001;
DRAM[54061] = 8'b11101001;
DRAM[54062] = 8'b11101010;
DRAM[54063] = 8'b11101011;
DRAM[54064] = 8'b11100101;
DRAM[54065] = 8'b11100100;
DRAM[54066] = 8'b11100010;
DRAM[54067] = 8'b11011111;
DRAM[54068] = 8'b11011100;
DRAM[54069] = 8'b11011001;
DRAM[54070] = 8'b11010111;
DRAM[54071] = 8'b11010101;
DRAM[54072] = 8'b11010010;
DRAM[54073] = 8'b11010001;
DRAM[54074] = 8'b11001001;
DRAM[54075] = 8'b11000001;
DRAM[54076] = 8'b11000001;
DRAM[54077] = 8'b11000111;
DRAM[54078] = 8'b11000110;
DRAM[54079] = 8'b10111111;
DRAM[54080] = 8'b10111100;
DRAM[54081] = 8'b10111110;
DRAM[54082] = 8'b10111010;
DRAM[54083] = 8'b10110000;
DRAM[54084] = 8'b10101011;
DRAM[54085] = 8'b10101111;
DRAM[54086] = 8'b10110100;
DRAM[54087] = 8'b10110100;
DRAM[54088] = 8'b10101101;
DRAM[54089] = 8'b10101100;
DRAM[54090] = 8'b10101000;
DRAM[54091] = 8'b10100110;
DRAM[54092] = 8'b10101000;
DRAM[54093] = 8'b10101100;
DRAM[54094] = 8'b10101000;
DRAM[54095] = 8'b10100001;
DRAM[54096] = 8'b10100000;
DRAM[54097] = 8'b10010110;
DRAM[54098] = 8'b10011001;
DRAM[54099] = 8'b10100001;
DRAM[54100] = 8'b10011101;
DRAM[54101] = 8'b10011010;
DRAM[54102] = 8'b10010110;
DRAM[54103] = 8'b10001101;
DRAM[54104] = 8'b10011001;
DRAM[54105] = 8'b10001001;
DRAM[54106] = 8'b10010010;
DRAM[54107] = 8'b10010010;
DRAM[54108] = 8'b1111010;
DRAM[54109] = 8'b1111110;
DRAM[54110] = 8'b10001100;
DRAM[54111] = 8'b10000000;
DRAM[54112] = 8'b1110000;
DRAM[54113] = 8'b1110000;
DRAM[54114] = 8'b1110110;
DRAM[54115] = 8'b1100110;
DRAM[54116] = 8'b1101001;
DRAM[54117] = 8'b1111111;
DRAM[54118] = 8'b1111101;
DRAM[54119] = 8'b1111101;
DRAM[54120] = 8'b1110011;
DRAM[54121] = 8'b1111000;
DRAM[54122] = 8'b1101110;
DRAM[54123] = 8'b1100100;
DRAM[54124] = 8'b1101001;
DRAM[54125] = 8'b1101100;
DRAM[54126] = 8'b1100111;
DRAM[54127] = 8'b1100101;
DRAM[54128] = 8'b1011001;
DRAM[54129] = 8'b1100101;
DRAM[54130] = 8'b1100010;
DRAM[54131] = 8'b1011010;
DRAM[54132] = 8'b1100001;
DRAM[54133] = 8'b1011111;
DRAM[54134] = 8'b1100100;
DRAM[54135] = 8'b1101000;
DRAM[54136] = 8'b1101000;
DRAM[54137] = 8'b1100001;
DRAM[54138] = 8'b1011010;
DRAM[54139] = 8'b1011011;
DRAM[54140] = 8'b1100001;
DRAM[54141] = 8'b1100010;
DRAM[54142] = 8'b1011001;
DRAM[54143] = 8'b1001110;
DRAM[54144] = 8'b1011010;
DRAM[54145] = 8'b1011100;
DRAM[54146] = 8'b1100101;
DRAM[54147] = 8'b1100110;
DRAM[54148] = 8'b1011111;
DRAM[54149] = 8'b1100011;
DRAM[54150] = 8'b1101000;
DRAM[54151] = 8'b1100000;
DRAM[54152] = 8'b1011010;
DRAM[54153] = 8'b1011101;
DRAM[54154] = 8'b1100100;
DRAM[54155] = 8'b1100100;
DRAM[54156] = 8'b1011111;
DRAM[54157] = 8'b1100111;
DRAM[54158] = 8'b1101100;
DRAM[54159] = 8'b1100011;
DRAM[54160] = 8'b1110000;
DRAM[54161] = 8'b1101001;
DRAM[54162] = 8'b1100010;
DRAM[54163] = 8'b1100010;
DRAM[54164] = 8'b1101001;
DRAM[54165] = 8'b1110010;
DRAM[54166] = 8'b1110101;
DRAM[54167] = 8'b1110100;
DRAM[54168] = 8'b1101011;
DRAM[54169] = 8'b1111010;
DRAM[54170] = 8'b1111100;
DRAM[54171] = 8'b10000001;
DRAM[54172] = 8'b1110011;
DRAM[54173] = 8'b1111011;
DRAM[54174] = 8'b1111000;
DRAM[54175] = 8'b1111011;
DRAM[54176] = 8'b1111110;
DRAM[54177] = 8'b10000000;
DRAM[54178] = 8'b10000010;
DRAM[54179] = 8'b10000011;
DRAM[54180] = 8'b10000011;
DRAM[54181] = 8'b10000101;
DRAM[54182] = 8'b10000111;
DRAM[54183] = 8'b10001010;
DRAM[54184] = 8'b10010101;
DRAM[54185] = 8'b10011110;
DRAM[54186] = 8'b10011111;
DRAM[54187] = 8'b10100100;
DRAM[54188] = 8'b10110000;
DRAM[54189] = 8'b10110011;
DRAM[54190] = 8'b10110011;
DRAM[54191] = 8'b10111010;
DRAM[54192] = 8'b10111011;
DRAM[54193] = 8'b10111010;
DRAM[54194] = 8'b10111100;
DRAM[54195] = 8'b11000010;
DRAM[54196] = 8'b11001011;
DRAM[54197] = 8'b11010001;
DRAM[54198] = 8'b11010011;
DRAM[54199] = 8'b11010011;
DRAM[54200] = 8'b11010111;
DRAM[54201] = 8'b11011010;
DRAM[54202] = 8'b11011110;
DRAM[54203] = 8'b11100010;
DRAM[54204] = 8'b11100110;
DRAM[54205] = 8'b11101010;
DRAM[54206] = 8'b11101101;
DRAM[54207] = 8'b11101111;
DRAM[54208] = 8'b11101101;
DRAM[54209] = 8'b11101001;
DRAM[54210] = 8'b11100000;
DRAM[54211] = 8'b11010001;
DRAM[54212] = 8'b11000000;
DRAM[54213] = 8'b10110000;
DRAM[54214] = 8'b10100010;
DRAM[54215] = 8'b10011001;
DRAM[54216] = 8'b10000111;
DRAM[54217] = 8'b10000101;
DRAM[54218] = 8'b10000010;
DRAM[54219] = 8'b1111111;
DRAM[54220] = 8'b1111101;
DRAM[54221] = 8'b1111100;
DRAM[54222] = 8'b1111101;
DRAM[54223] = 8'b1111111;
DRAM[54224] = 8'b1111000;
DRAM[54225] = 8'b1111010;
DRAM[54226] = 8'b1111001;
DRAM[54227] = 8'b1110101;
DRAM[54228] = 8'b1110101;
DRAM[54229] = 8'b1111000;
DRAM[54230] = 8'b1111001;
DRAM[54231] = 8'b1110110;
DRAM[54232] = 8'b1110100;
DRAM[54233] = 8'b1110011;
DRAM[54234] = 8'b1110001;
DRAM[54235] = 8'b1110000;
DRAM[54236] = 8'b1101111;
DRAM[54237] = 8'b1101111;
DRAM[54238] = 8'b1110000;
DRAM[54239] = 8'b1110001;
DRAM[54240] = 8'b1110010;
DRAM[54241] = 8'b1110010;
DRAM[54242] = 8'b1110010;
DRAM[54243] = 8'b1110001;
DRAM[54244] = 8'b1110010;
DRAM[54245] = 8'b1110010;
DRAM[54246] = 8'b1110011;
DRAM[54247] = 8'b1110100;
DRAM[54248] = 8'b1110110;
DRAM[54249] = 8'b1110110;
DRAM[54250] = 8'b1110110;
DRAM[54251] = 8'b1110110;
DRAM[54252] = 8'b1110101;
DRAM[54253] = 8'b1110100;
DRAM[54254] = 8'b1110010;
DRAM[54255] = 8'b1110010;
DRAM[54256] = 8'b1110000;
DRAM[54257] = 8'b1110000;
DRAM[54258] = 8'b1110000;
DRAM[54259] = 8'b1110000;
DRAM[54260] = 8'b1101111;
DRAM[54261] = 8'b1101110;
DRAM[54262] = 8'b1101100;
DRAM[54263] = 8'b1101100;
DRAM[54264] = 8'b1101011;
DRAM[54265] = 8'b1101100;
DRAM[54266] = 8'b1101100;
DRAM[54267] = 8'b1101101;
DRAM[54268] = 8'b1101110;
DRAM[54269] = 8'b1101111;
DRAM[54270] = 8'b1101111;
DRAM[54271] = 8'b1101111;
DRAM[54272] = 8'b10011001;
DRAM[54273] = 8'b10011001;
DRAM[54274] = 8'b10011001;
DRAM[54275] = 8'b10011001;
DRAM[54276] = 8'b10011001;
DRAM[54277] = 8'b10011000;
DRAM[54278] = 8'b10011000;
DRAM[54279] = 8'b10011000;
DRAM[54280] = 8'b10011101;
DRAM[54281] = 8'b10011110;
DRAM[54282] = 8'b10011111;
DRAM[54283] = 8'b10011101;
DRAM[54284] = 8'b10011011;
DRAM[54285] = 8'b10011001;
DRAM[54286] = 8'b10011010;
DRAM[54287] = 8'b10011011;
DRAM[54288] = 8'b10011001;
DRAM[54289] = 8'b10011001;
DRAM[54290] = 8'b10011001;
DRAM[54291] = 8'b10011001;
DRAM[54292] = 8'b10100000;
DRAM[54293] = 8'b10110100;
DRAM[54294] = 8'b11010101;
DRAM[54295] = 8'b11110000;
DRAM[54296] = 8'b11111001;
DRAM[54297] = 8'b11111110;
DRAM[54298] = 8'b11111111;
DRAM[54299] = 8'b11111111;
DRAM[54300] = 8'b11111101;
DRAM[54301] = 8'b11111100;
DRAM[54302] = 8'b11111010;
DRAM[54303] = 8'b11110111;
DRAM[54304] = 8'b11111100;
DRAM[54305] = 8'b11111011;
DRAM[54306] = 8'b11111011;
DRAM[54307] = 8'b11111011;
DRAM[54308] = 8'b11111011;
DRAM[54309] = 8'b11111010;
DRAM[54310] = 8'b11110110;
DRAM[54311] = 8'b11110011;
DRAM[54312] = 8'b11100110;
DRAM[54313] = 8'b11100110;
DRAM[54314] = 8'b11100110;
DRAM[54315] = 8'b11100101;
DRAM[54316] = 8'b11100101;
DRAM[54317] = 8'b11100100;
DRAM[54318] = 8'b11100100;
DRAM[54319] = 8'b11100011;
DRAM[54320] = 8'b11100111;
DRAM[54321] = 8'b11100101;
DRAM[54322] = 8'b11100010;
DRAM[54323] = 8'b11011110;
DRAM[54324] = 8'b11011001;
DRAM[54325] = 8'b11010101;
DRAM[54326] = 8'b11010001;
DRAM[54327] = 8'b11001111;
DRAM[54328] = 8'b11001100;
DRAM[54329] = 8'b11000001;
DRAM[54330] = 8'b10111011;
DRAM[54331] = 8'b10111101;
DRAM[54332] = 8'b10111111;
DRAM[54333] = 8'b10111011;
DRAM[54334] = 8'b10111011;
DRAM[54335] = 8'b10111110;
DRAM[54336] = 8'b10111111;
DRAM[54337] = 8'b10111110;
DRAM[54338] = 8'b10111000;
DRAM[54339] = 8'b10101110;
DRAM[54340] = 8'b10101001;
DRAM[54341] = 8'b10101010;
DRAM[54342] = 8'b10101011;
DRAM[54343] = 8'b10101011;
DRAM[54344] = 8'b10101101;
DRAM[54345] = 8'b10011111;
DRAM[54346] = 8'b10011101;
DRAM[54347] = 8'b10101100;
DRAM[54348] = 8'b10110100;
DRAM[54349] = 8'b10101100;
DRAM[54350] = 8'b10100010;
DRAM[54351] = 8'b10100000;
DRAM[54352] = 8'b10011111;
DRAM[54353] = 8'b10010111;
DRAM[54354] = 8'b10011100;
DRAM[54355] = 8'b10011111;
DRAM[54356] = 8'b10010101;
DRAM[54357] = 8'b10010000;
DRAM[54358] = 8'b10010001;
DRAM[54359] = 8'b10001101;
DRAM[54360] = 8'b10011010;
DRAM[54361] = 8'b10001000;
DRAM[54362] = 8'b10010000;
DRAM[54363] = 8'b10010011;
DRAM[54364] = 8'b1111101;
DRAM[54365] = 8'b10000000;
DRAM[54366] = 8'b10001000;
DRAM[54367] = 8'b1110111;
DRAM[54368] = 8'b1110011;
DRAM[54369] = 8'b1110100;
DRAM[54370] = 8'b1111010;
DRAM[54371] = 8'b1101010;
DRAM[54372] = 8'b1101011;
DRAM[54373] = 8'b10000000;
DRAM[54374] = 8'b1111111;
DRAM[54375] = 8'b10000000;
DRAM[54376] = 8'b1110101;
DRAM[54377] = 8'b1110011;
DRAM[54378] = 8'b1100111;
DRAM[54379] = 8'b1011111;
DRAM[54380] = 8'b1100110;
DRAM[54381] = 8'b1101000;
DRAM[54382] = 8'b1100101;
DRAM[54383] = 8'b1100111;
DRAM[54384] = 8'b1010111;
DRAM[54385] = 8'b1100000;
DRAM[54386] = 8'b1011101;
DRAM[54387] = 8'b1011001;
DRAM[54388] = 8'b1011111;
DRAM[54389] = 8'b1100111;
DRAM[54390] = 8'b1100001;
DRAM[54391] = 8'b1101000;
DRAM[54392] = 8'b1100100;
DRAM[54393] = 8'b1011111;
DRAM[54394] = 8'b1011011;
DRAM[54395] = 8'b1011100;
DRAM[54396] = 8'b1011110;
DRAM[54397] = 8'b1011101;
DRAM[54398] = 8'b1011000;
DRAM[54399] = 8'b1010101;
DRAM[54400] = 8'b1011011;
DRAM[54401] = 8'b1011100;
DRAM[54402] = 8'b1100110;
DRAM[54403] = 8'b1101000;
DRAM[54404] = 8'b1100011;
DRAM[54405] = 8'b1100111;
DRAM[54406] = 8'b1101010;
DRAM[54407] = 8'b1100000;
DRAM[54408] = 8'b1100011;
DRAM[54409] = 8'b1010111;
DRAM[54410] = 8'b1011100;
DRAM[54411] = 8'b1101000;
DRAM[54412] = 8'b1101001;
DRAM[54413] = 8'b1101001;
DRAM[54414] = 8'b1101010;
DRAM[54415] = 8'b1100101;
DRAM[54416] = 8'b1101100;
DRAM[54417] = 8'b1101001;
DRAM[54418] = 8'b1100110;
DRAM[54419] = 8'b1100110;
DRAM[54420] = 8'b1101000;
DRAM[54421] = 8'b1101101;
DRAM[54422] = 8'b1110100;
DRAM[54423] = 8'b1111010;
DRAM[54424] = 8'b1101011;
DRAM[54425] = 8'b1101111;
DRAM[54426] = 8'b1111011;
DRAM[54427] = 8'b1110100;
DRAM[54428] = 8'b1111110;
DRAM[54429] = 8'b1111010;
DRAM[54430] = 8'b10000100;
DRAM[54431] = 8'b10000010;
DRAM[54432] = 8'b10000001;
DRAM[54433] = 8'b10000011;
DRAM[54434] = 8'b10000101;
DRAM[54435] = 8'b10000110;
DRAM[54436] = 8'b10000110;
DRAM[54437] = 8'b10000111;
DRAM[54438] = 8'b10001001;
DRAM[54439] = 8'b10001011;
DRAM[54440] = 8'b10001011;
DRAM[54441] = 8'b10010010;
DRAM[54442] = 8'b10010010;
DRAM[54443] = 8'b10010111;
DRAM[54444] = 8'b10100110;
DRAM[54445] = 8'b10101110;
DRAM[54446] = 8'b10110011;
DRAM[54447] = 8'b10111110;
DRAM[54448] = 8'b10111101;
DRAM[54449] = 8'b10111100;
DRAM[54450] = 8'b10111101;
DRAM[54451] = 8'b11000011;
DRAM[54452] = 8'b11001011;
DRAM[54453] = 8'b11010001;
DRAM[54454] = 8'b11010011;
DRAM[54455] = 8'b11010010;
DRAM[54456] = 8'b11010101;
DRAM[54457] = 8'b11010100;
DRAM[54458] = 8'b11010101;
DRAM[54459] = 8'b11011100;
DRAM[54460] = 8'b11100110;
DRAM[54461] = 8'b11101110;
DRAM[54462] = 8'b11110000;
DRAM[54463] = 8'b11101111;
DRAM[54464] = 8'b11110001;
DRAM[54465] = 8'b11011000;
DRAM[54466] = 8'b10111111;
DRAM[54467] = 8'b10111100;
DRAM[54468] = 8'b11000101;
DRAM[54469] = 8'b11000111;
DRAM[54470] = 8'b10110111;
DRAM[54471] = 8'b10100110;
DRAM[54472] = 8'b10011000;
DRAM[54473] = 8'b10010000;
DRAM[54474] = 8'b10000110;
DRAM[54475] = 8'b10000001;
DRAM[54476] = 8'b10000000;
DRAM[54477] = 8'b1111111;
DRAM[54478] = 8'b1111100;
DRAM[54479] = 8'b1111001;
DRAM[54480] = 8'b1111001;
DRAM[54481] = 8'b1111011;
DRAM[54482] = 8'b1111010;
DRAM[54483] = 8'b1110110;
DRAM[54484] = 8'b1110110;
DRAM[54485] = 8'b1111001;
DRAM[54486] = 8'b1111001;
DRAM[54487] = 8'b1110111;
DRAM[54488] = 8'b1110101;
DRAM[54489] = 8'b1110100;
DRAM[54490] = 8'b1110010;
DRAM[54491] = 8'b1110000;
DRAM[54492] = 8'b1101111;
DRAM[54493] = 8'b1101111;
DRAM[54494] = 8'b1110000;
DRAM[54495] = 8'b1110000;
DRAM[54496] = 8'b1110001;
DRAM[54497] = 8'b1110001;
DRAM[54498] = 8'b1110000;
DRAM[54499] = 8'b1110001;
DRAM[54500] = 8'b1110001;
DRAM[54501] = 8'b1110010;
DRAM[54502] = 8'b1110011;
DRAM[54503] = 8'b1110100;
DRAM[54504] = 8'b1110101;
DRAM[54505] = 8'b1110101;
DRAM[54506] = 8'b1110101;
DRAM[54507] = 8'b1110101;
DRAM[54508] = 8'b1110100;
DRAM[54509] = 8'b1110011;
DRAM[54510] = 8'b1110010;
DRAM[54511] = 8'b1110001;
DRAM[54512] = 8'b1101111;
DRAM[54513] = 8'b1101111;
DRAM[54514] = 8'b1101111;
DRAM[54515] = 8'b1101111;
DRAM[54516] = 8'b1101110;
DRAM[54517] = 8'b1101101;
DRAM[54518] = 8'b1101011;
DRAM[54519] = 8'b1101011;
DRAM[54520] = 8'b1101011;
DRAM[54521] = 8'b1101011;
DRAM[54522] = 8'b1101011;
DRAM[54523] = 8'b1101100;
DRAM[54524] = 8'b1101101;
DRAM[54525] = 8'b1101110;
DRAM[54526] = 8'b1101110;
DRAM[54527] = 8'b1101111;
DRAM[54528] = 8'b10011001;
DRAM[54529] = 8'b10011001;
DRAM[54530] = 8'b10011010;
DRAM[54531] = 8'b10011010;
DRAM[54532] = 8'b10011010;
DRAM[54533] = 8'b10011010;
DRAM[54534] = 8'b10011010;
DRAM[54535] = 8'b10011010;
DRAM[54536] = 8'b10011110;
DRAM[54537] = 8'b10011111;
DRAM[54538] = 8'b10011111;
DRAM[54539] = 8'b10011110;
DRAM[54540] = 8'b10011100;
DRAM[54541] = 8'b10011010;
DRAM[54542] = 8'b10011011;
DRAM[54543] = 8'b10011100;
DRAM[54544] = 8'b10010110;
DRAM[54545] = 8'b10010111;
DRAM[54546] = 8'b10011010;
DRAM[54547] = 8'b10100001;
DRAM[54548] = 8'b10110000;
DRAM[54549] = 8'b11001001;
DRAM[54550] = 8'b11101000;
DRAM[54551] = 8'b11111101;
DRAM[54552] = 8'b11111000;
DRAM[54553] = 8'b11111100;
DRAM[54554] = 8'b11111111;
DRAM[54555] = 8'b11111111;
DRAM[54556] = 8'b11111101;
DRAM[54557] = 8'b11111010;
DRAM[54558] = 8'b11111001;
DRAM[54559] = 8'b11111001;
DRAM[54560] = 8'b11111100;
DRAM[54561] = 8'b11111010;
DRAM[54562] = 8'b11110111;
DRAM[54563] = 8'b11110101;
DRAM[54564] = 8'b11110011;
DRAM[54565] = 8'b11110001;
DRAM[54566] = 8'b11101101;
DRAM[54567] = 8'b11101001;
DRAM[54568] = 8'b11100100;
DRAM[54569] = 8'b11100100;
DRAM[54570] = 8'b11100100;
DRAM[54571] = 8'b11100100;
DRAM[54572] = 8'b11100011;
DRAM[54573] = 8'b11100010;
DRAM[54574] = 8'b11100001;
DRAM[54575] = 8'b11100001;
DRAM[54576] = 8'b11100101;
DRAM[54577] = 8'b11100011;
DRAM[54578] = 8'b11011111;
DRAM[54579] = 8'b11011010;
DRAM[54580] = 8'b11010101;
DRAM[54581] = 8'b11010000;
DRAM[54582] = 8'b11001100;
DRAM[54583] = 8'b11001010;
DRAM[54584] = 8'b11000110;
DRAM[54585] = 8'b10110101;
DRAM[54586] = 8'b10101011;
DRAM[54587] = 8'b10101111;
DRAM[54588] = 8'b10101111;
DRAM[54589] = 8'b10101001;
DRAM[54590] = 8'b10101011;
DRAM[54591] = 8'b10110100;
DRAM[54592] = 8'b10110000;
DRAM[54593] = 8'b10101101;
DRAM[54594] = 8'b10101000;
DRAM[54595] = 8'b10100010;
DRAM[54596] = 8'b10011101;
DRAM[54597] = 8'b10011100;
DRAM[54598] = 8'b10011011;
DRAM[54599] = 8'b10011011;
DRAM[54600] = 8'b10101110;
DRAM[54601] = 8'b10011010;
DRAM[54602] = 8'b10010110;
DRAM[54603] = 8'b10101000;
DRAM[54604] = 8'b10101111;
DRAM[54605] = 8'b10100010;
DRAM[54606] = 8'b10011101;
DRAM[54607] = 8'b10100101;
DRAM[54608] = 8'b10100101;
DRAM[54609] = 8'b10011011;
DRAM[54610] = 8'b10011010;
DRAM[54611] = 8'b10011001;
DRAM[54612] = 8'b10001110;
DRAM[54613] = 8'b10001101;
DRAM[54614] = 8'b10010110;
DRAM[54615] = 8'b10011000;
DRAM[54616] = 8'b10011000;
DRAM[54617] = 8'b10001100;
DRAM[54618] = 8'b10010000;
DRAM[54619] = 8'b10010000;
DRAM[54620] = 8'b10000010;
DRAM[54621] = 8'b10000001;
DRAM[54622] = 8'b10000100;
DRAM[54623] = 8'b1110111;
DRAM[54624] = 8'b1111001;
DRAM[54625] = 8'b1110101;
DRAM[54626] = 8'b1111010;
DRAM[54627] = 8'b1101101;
DRAM[54628] = 8'b1101111;
DRAM[54629] = 8'b1111111;
DRAM[54630] = 8'b1111101;
DRAM[54631] = 8'b10000001;
DRAM[54632] = 8'b1110110;
DRAM[54633] = 8'b1101010;
DRAM[54634] = 8'b1100010;
DRAM[54635] = 8'b1100000;
DRAM[54636] = 8'b1100001;
DRAM[54637] = 8'b1100001;
DRAM[54638] = 8'b1100000;
DRAM[54639] = 8'b1011111;
DRAM[54640] = 8'b1011011;
DRAM[54641] = 8'b1011100;
DRAM[54642] = 8'b1011000;
DRAM[54643] = 8'b1011010;
DRAM[54644] = 8'b1011101;
DRAM[54645] = 8'b1101010;
DRAM[54646] = 8'b1011000;
DRAM[54647] = 8'b1100101;
DRAM[54648] = 8'b1100101;
DRAM[54649] = 8'b1100001;
DRAM[54650] = 8'b1011110;
DRAM[54651] = 8'b1011111;
DRAM[54652] = 8'b1011110;
DRAM[54653] = 8'b1011010;
DRAM[54654] = 8'b1011010;
DRAM[54655] = 8'b1011100;
DRAM[54656] = 8'b1011010;
DRAM[54657] = 8'b1011011;
DRAM[54658] = 8'b1100100;
DRAM[54659] = 8'b1100111;
DRAM[54660] = 8'b1100011;
DRAM[54661] = 8'b1101000;
DRAM[54662] = 8'b1101011;
DRAM[54663] = 8'b1100001;
DRAM[54664] = 8'b1100111;
DRAM[54665] = 8'b1010011;
DRAM[54666] = 8'b1010011;
DRAM[54667] = 8'b1100011;
DRAM[54668] = 8'b1100110;
DRAM[54669] = 8'b1100101;
DRAM[54670] = 8'b1100110;
DRAM[54671] = 8'b1100100;
DRAM[54672] = 8'b1011110;
DRAM[54673] = 8'b1100111;
DRAM[54674] = 8'b1110000;
DRAM[54675] = 8'b1101111;
DRAM[54676] = 8'b1100101;
DRAM[54677] = 8'b1100010;
DRAM[54678] = 8'b1101110;
DRAM[54679] = 8'b1111111;
DRAM[54680] = 8'b10000010;
DRAM[54681] = 8'b1111001;
DRAM[54682] = 8'b1111110;
DRAM[54683] = 8'b1101101;
DRAM[54684] = 8'b1111011;
DRAM[54685] = 8'b1110010;
DRAM[54686] = 8'b10000010;
DRAM[54687] = 8'b10000000;
DRAM[54688] = 8'b10000101;
DRAM[54689] = 8'b10001000;
DRAM[54690] = 8'b10001100;
DRAM[54691] = 8'b10001110;
DRAM[54692] = 8'b10001111;
DRAM[54693] = 8'b10010001;
DRAM[54694] = 8'b10010011;
DRAM[54695] = 8'b10010101;
DRAM[54696] = 8'b10001100;
DRAM[54697] = 8'b10010001;
DRAM[54698] = 8'b10001110;
DRAM[54699] = 8'b10001111;
DRAM[54700] = 8'b10011011;
DRAM[54701] = 8'b10100010;
DRAM[54702] = 8'b10100111;
DRAM[54703] = 8'b10110010;
DRAM[54704] = 8'b10111010;
DRAM[54705] = 8'b10111011;
DRAM[54706] = 8'b10111111;
DRAM[54707] = 8'b11000101;
DRAM[54708] = 8'b11001100;
DRAM[54709] = 8'b11010010;
DRAM[54710] = 8'b11010101;
DRAM[54711] = 8'b11010110;
DRAM[54712] = 8'b11011011;
DRAM[54713] = 8'b11011000;
DRAM[54714] = 8'b11011000;
DRAM[54715] = 8'b11011101;
DRAM[54716] = 8'b11100111;
DRAM[54717] = 8'b11101110;
DRAM[54718] = 8'b11110001;
DRAM[54719] = 8'b11110001;
DRAM[54720] = 8'b11111111;
DRAM[54721] = 8'b11011111;
DRAM[54722] = 8'b10111100;
DRAM[54723] = 8'b10101100;
DRAM[54724] = 8'b10101100;
DRAM[54725] = 8'b10101110;
DRAM[54726] = 8'b10101100;
DRAM[54727] = 8'b10101001;
DRAM[54728] = 8'b10100001;
DRAM[54729] = 8'b10010111;
DRAM[54730] = 8'b10001100;
DRAM[54731] = 8'b10000110;
DRAM[54732] = 8'b10000110;
DRAM[54733] = 8'b10000101;
DRAM[54734] = 8'b10000000;
DRAM[54735] = 8'b1111011;
DRAM[54736] = 8'b1111010;
DRAM[54737] = 8'b1111100;
DRAM[54738] = 8'b1111011;
DRAM[54739] = 8'b1110111;
DRAM[54740] = 8'b1110111;
DRAM[54741] = 8'b1111010;
DRAM[54742] = 8'b1111010;
DRAM[54743] = 8'b1110111;
DRAM[54744] = 8'b1110110;
DRAM[54745] = 8'b1110101;
DRAM[54746] = 8'b1110011;
DRAM[54747] = 8'b1110001;
DRAM[54748] = 8'b1101111;
DRAM[54749] = 8'b1101111;
DRAM[54750] = 8'b1110000;
DRAM[54751] = 8'b1110000;
DRAM[54752] = 8'b1110000;
DRAM[54753] = 8'b1110000;
DRAM[54754] = 8'b1101111;
DRAM[54755] = 8'b1110000;
DRAM[54756] = 8'b1110000;
DRAM[54757] = 8'b1110010;
DRAM[54758] = 8'b1110011;
DRAM[54759] = 8'b1110011;
DRAM[54760] = 8'b1110100;
DRAM[54761] = 8'b1110100;
DRAM[54762] = 8'b1110100;
DRAM[54763] = 8'b1110100;
DRAM[54764] = 8'b1110011;
DRAM[54765] = 8'b1110001;
DRAM[54766] = 8'b1110000;
DRAM[54767] = 8'b1101111;
DRAM[54768] = 8'b1101110;
DRAM[54769] = 8'b1101110;
DRAM[54770] = 8'b1101110;
DRAM[54771] = 8'b1101110;
DRAM[54772] = 8'b1101101;
DRAM[54773] = 8'b1101100;
DRAM[54774] = 8'b1101011;
DRAM[54775] = 8'b1101010;
DRAM[54776] = 8'b1101010;
DRAM[54777] = 8'b1101010;
DRAM[54778] = 8'b1101011;
DRAM[54779] = 8'b1101011;
DRAM[54780] = 8'b1101100;
DRAM[54781] = 8'b1101101;
DRAM[54782] = 8'b1101110;
DRAM[54783] = 8'b1101110;
DRAM[54784] = 8'b10011001;
DRAM[54785] = 8'b10011001;
DRAM[54786] = 8'b10011010;
DRAM[54787] = 8'b10011010;
DRAM[54788] = 8'b10011011;
DRAM[54789] = 8'b10011100;
DRAM[54790] = 8'b10011100;
DRAM[54791] = 8'b10011100;
DRAM[54792] = 8'b10011110;
DRAM[54793] = 8'b10011111;
DRAM[54794] = 8'b10100000;
DRAM[54795] = 8'b10011110;
DRAM[54796] = 8'b10011100;
DRAM[54797] = 8'b10011010;
DRAM[54798] = 8'b10011011;
DRAM[54799] = 8'b10011100;
DRAM[54800] = 8'b10010111;
DRAM[54801] = 8'b10011010;
DRAM[54802] = 8'b10100001;
DRAM[54803] = 8'b10101111;
DRAM[54804] = 8'b11000110;
DRAM[54805] = 8'b11100000;
DRAM[54806] = 8'b11110100;
DRAM[54807] = 8'b11111110;
DRAM[54808] = 8'b11111100;
DRAM[54809] = 8'b11111100;
DRAM[54810] = 8'b11111101;
DRAM[54811] = 8'b11111110;
DRAM[54812] = 8'b11111100;
DRAM[54813] = 8'b11111010;
DRAM[54814] = 8'b11111001;
DRAM[54815] = 8'b11111001;
DRAM[54816] = 8'b11111100;
DRAM[54817] = 8'b11111001;
DRAM[54818] = 8'b11110100;
DRAM[54819] = 8'b11101111;
DRAM[54820] = 8'b11101100;
DRAM[54821] = 8'b11101000;
DRAM[54822] = 8'b11100100;
DRAM[54823] = 8'b11100001;
DRAM[54824] = 8'b11101011;
DRAM[54825] = 8'b11101001;
DRAM[54826] = 8'b11100111;
DRAM[54827] = 8'b11100101;
DRAM[54828] = 8'b11100100;
DRAM[54829] = 8'b11100100;
DRAM[54830] = 8'b11100101;
DRAM[54831] = 8'b11100110;
DRAM[54832] = 8'b11011110;
DRAM[54833] = 8'b11011100;
DRAM[54834] = 8'b11011001;
DRAM[54835] = 8'b11010101;
DRAM[54836] = 8'b11010000;
DRAM[54837] = 8'b11001100;
DRAM[54838] = 8'b11001000;
DRAM[54839] = 8'b11000111;
DRAM[54840] = 8'b11000000;
DRAM[54841] = 8'b10111000;
DRAM[54842] = 8'b10110010;
DRAM[54843] = 8'b10110001;
DRAM[54844] = 8'b10110001;
DRAM[54845] = 8'b10101111;
DRAM[54846] = 8'b10101101;
DRAM[54847] = 8'b10101101;
DRAM[54848] = 8'b10101000;
DRAM[54849] = 8'b10100110;
DRAM[54850] = 8'b10100100;
DRAM[54851] = 8'b10100101;
DRAM[54852] = 8'b10100101;
DRAM[54853] = 8'b10100110;
DRAM[54854] = 8'b10100110;
DRAM[54855] = 8'b10100111;
DRAM[54856] = 8'b10100101;
DRAM[54857] = 8'b10011110;
DRAM[54858] = 8'b10011111;
DRAM[54859] = 8'b10100110;
DRAM[54860] = 8'b10100100;
DRAM[54861] = 8'b10011001;
DRAM[54862] = 8'b10011001;
DRAM[54863] = 8'b10100011;
DRAM[54864] = 8'b10100001;
DRAM[54865] = 8'b10010110;
DRAM[54866] = 8'b10010110;
DRAM[54867] = 8'b10011001;
DRAM[54868] = 8'b10010100;
DRAM[54869] = 8'b10010111;
DRAM[54870] = 8'b10011111;
DRAM[54871] = 8'b10011110;
DRAM[54872] = 8'b10010100;
DRAM[54873] = 8'b10010100;
DRAM[54874] = 8'b10010011;
DRAM[54875] = 8'b10001101;
DRAM[54876] = 8'b10000101;
DRAM[54877] = 8'b10000001;
DRAM[54878] = 8'b10000010;
DRAM[54879] = 8'b10000010;
DRAM[54880] = 8'b1111111;
DRAM[54881] = 8'b1110100;
DRAM[54882] = 8'b1110111;
DRAM[54883] = 8'b1101111;
DRAM[54884] = 8'b1110010;
DRAM[54885] = 8'b1111101;
DRAM[54886] = 8'b1111001;
DRAM[54887] = 8'b10000000;
DRAM[54888] = 8'b1111010;
DRAM[54889] = 8'b1100101;
DRAM[54890] = 8'b1100101;
DRAM[54891] = 8'b1101011;
DRAM[54892] = 8'b1100001;
DRAM[54893] = 8'b1011110;
DRAM[54894] = 8'b1011110;
DRAM[54895] = 8'b1010001;
DRAM[54896] = 8'b1100000;
DRAM[54897] = 8'b1011010;
DRAM[54898] = 8'b1011000;
DRAM[54899] = 8'b1011110;
DRAM[54900] = 8'b1011001;
DRAM[54901] = 8'b1100100;
DRAM[54902] = 8'b1001011;
DRAM[54903] = 8'b1100001;
DRAM[54904] = 8'b1101010;
DRAM[54905] = 8'b1100100;
DRAM[54906] = 8'b1100000;
DRAM[54907] = 8'b1100010;
DRAM[54908] = 8'b1100001;
DRAM[54909] = 8'b1011101;
DRAM[54910] = 8'b1011101;
DRAM[54911] = 8'b1100000;
DRAM[54912] = 8'b1010111;
DRAM[54913] = 8'b1010111;
DRAM[54914] = 8'b1011111;
DRAM[54915] = 8'b1100011;
DRAM[54916] = 8'b1100001;
DRAM[54917] = 8'b1100111;
DRAM[54918] = 8'b1101010;
DRAM[54919] = 8'b1100000;
DRAM[54920] = 8'b1100110;
DRAM[54921] = 8'b1010111;
DRAM[54922] = 8'b1010100;
DRAM[54923] = 8'b1010111;
DRAM[54924] = 8'b1011000;
DRAM[54925] = 8'b1100000;
DRAM[54926] = 8'b1101000;
DRAM[54927] = 8'b1100100;
DRAM[54928] = 8'b1011010;
DRAM[54929] = 8'b1011111;
DRAM[54930] = 8'b1101001;
DRAM[54931] = 8'b1101110;
DRAM[54932] = 8'b1101010;
DRAM[54933] = 8'b1100100;
DRAM[54934] = 8'b1101010;
DRAM[54935] = 8'b1110100;
DRAM[54936] = 8'b10000101;
DRAM[54937] = 8'b10000001;
DRAM[54938] = 8'b1111111;
DRAM[54939] = 8'b1111000;
DRAM[54940] = 8'b1111000;
DRAM[54941] = 8'b1110101;
DRAM[54942] = 8'b1111100;
DRAM[54943] = 8'b10000000;
DRAM[54944] = 8'b1111101;
DRAM[54945] = 8'b10000000;
DRAM[54946] = 8'b10000100;
DRAM[54947] = 8'b10000111;
DRAM[54948] = 8'b10000111;
DRAM[54949] = 8'b10001000;
DRAM[54950] = 8'b10001010;
DRAM[54951] = 8'b10001011;
DRAM[54952] = 8'b10010100;
DRAM[54953] = 8'b10011000;
DRAM[54954] = 8'b10010011;
DRAM[54955] = 8'b10010000;
DRAM[54956] = 8'b10011001;
DRAM[54957] = 8'b10011011;
DRAM[54958] = 8'b10011100;
DRAM[54959] = 8'b10100101;
DRAM[54960] = 8'b10101111;
DRAM[54961] = 8'b10110011;
DRAM[54962] = 8'b10111010;
DRAM[54963] = 8'b11000000;
DRAM[54964] = 8'b11000111;
DRAM[54965] = 8'b11001110;
DRAM[54966] = 8'b11010100;
DRAM[54967] = 8'b11011001;
DRAM[54968] = 8'b11011011;
DRAM[54969] = 8'b11011101;
DRAM[54970] = 8'b11100000;
DRAM[54971] = 8'b11100010;
DRAM[54972] = 8'b11100101;
DRAM[54973] = 8'b11101010;
DRAM[54974] = 8'b11110001;
DRAM[54975] = 8'b11110110;
DRAM[54976] = 8'b11111011;
DRAM[54977] = 8'b11101011;
DRAM[54978] = 8'b11010110;
DRAM[54979] = 8'b11000001;
DRAM[54980] = 8'b10101100;
DRAM[54981] = 8'b10011111;
DRAM[54982] = 8'b10011110;
DRAM[54983] = 8'b10100110;
DRAM[54984] = 8'b10010111;
DRAM[54985] = 8'b10010010;
DRAM[54986] = 8'b10001101;
DRAM[54987] = 8'b10001010;
DRAM[54988] = 8'b10001001;
DRAM[54989] = 8'b10000111;
DRAM[54990] = 8'b10000100;
DRAM[54991] = 8'b10000001;
DRAM[54992] = 8'b1111010;
DRAM[54993] = 8'b1111100;
DRAM[54994] = 8'b1111100;
DRAM[54995] = 8'b1111000;
DRAM[54996] = 8'b1110111;
DRAM[54997] = 8'b1111010;
DRAM[54998] = 8'b1111011;
DRAM[54999] = 8'b1111000;
DRAM[55000] = 8'b1110111;
DRAM[55001] = 8'b1110101;
DRAM[55002] = 8'b1110011;
DRAM[55003] = 8'b1110001;
DRAM[55004] = 8'b1110000;
DRAM[55005] = 8'b1101111;
DRAM[55006] = 8'b1110000;
DRAM[55007] = 8'b1110000;
DRAM[55008] = 8'b1101111;
DRAM[55009] = 8'b1101111;
DRAM[55010] = 8'b1101111;
DRAM[55011] = 8'b1101111;
DRAM[55012] = 8'b1110000;
DRAM[55013] = 8'b1110001;
DRAM[55014] = 8'b1110010;
DRAM[55015] = 8'b1110011;
DRAM[55016] = 8'b1110010;
DRAM[55017] = 8'b1110010;
DRAM[55018] = 8'b1110010;
DRAM[55019] = 8'b1110010;
DRAM[55020] = 8'b1110001;
DRAM[55021] = 8'b1110000;
DRAM[55022] = 8'b1101111;
DRAM[55023] = 8'b1101110;
DRAM[55024] = 8'b1101110;
DRAM[55025] = 8'b1101110;
DRAM[55026] = 8'b1101110;
DRAM[55027] = 8'b1101101;
DRAM[55028] = 8'b1101101;
DRAM[55029] = 8'b1101011;
DRAM[55030] = 8'b1101010;
DRAM[55031] = 8'b1101001;
DRAM[55032] = 8'b1101001;
DRAM[55033] = 8'b1101001;
DRAM[55034] = 8'b1101010;
DRAM[55035] = 8'b1101011;
DRAM[55036] = 8'b1101100;
DRAM[55037] = 8'b1101100;
DRAM[55038] = 8'b1101101;
DRAM[55039] = 8'b1101101;
DRAM[55040] = 8'b10011000;
DRAM[55041] = 8'b10011001;
DRAM[55042] = 8'b10011010;
DRAM[55043] = 8'b10011011;
DRAM[55044] = 8'b10011100;
DRAM[55045] = 8'b10011101;
DRAM[55046] = 8'b10011101;
DRAM[55047] = 8'b10011110;
DRAM[55048] = 8'b10011110;
DRAM[55049] = 8'b10011111;
DRAM[55050] = 8'b10100000;
DRAM[55051] = 8'b10011110;
DRAM[55052] = 8'b10011100;
DRAM[55053] = 8'b10011010;
DRAM[55054] = 8'b10011011;
DRAM[55055] = 8'b10011100;
DRAM[55056] = 8'b10011010;
DRAM[55057] = 8'b10011101;
DRAM[55058] = 8'b10100111;
DRAM[55059] = 8'b10111010;
DRAM[55060] = 8'b11010101;
DRAM[55061] = 8'b11101100;
DRAM[55062] = 8'b11110111;
DRAM[55063] = 8'b11111000;
DRAM[55064] = 8'b11111111;
DRAM[55065] = 8'b11111101;
DRAM[55066] = 8'b11111010;
DRAM[55067] = 8'b11111011;
DRAM[55068] = 8'b11111100;
DRAM[55069] = 8'b11111100;
DRAM[55070] = 8'b11111010;
DRAM[55071] = 8'b11111001;
DRAM[55072] = 8'b11111001;
DRAM[55073] = 8'b11110110;
DRAM[55074] = 8'b11110010;
DRAM[55075] = 8'b11110000;
DRAM[55076] = 8'b11110000;
DRAM[55077] = 8'b11110000;
DRAM[55078] = 8'b11110000;
DRAM[55079] = 8'b11101111;
DRAM[55080] = 8'b11101111;
DRAM[55081] = 8'b11101100;
DRAM[55082] = 8'b11100111;
DRAM[55083] = 8'b11100011;
DRAM[55084] = 8'b11100010;
DRAM[55085] = 8'b11100011;
DRAM[55086] = 8'b11100110;
DRAM[55087] = 8'b11101000;
DRAM[55088] = 8'b11011000;
DRAM[55089] = 8'b11010110;
DRAM[55090] = 8'b11010100;
DRAM[55091] = 8'b11010000;
DRAM[55092] = 8'b11001101;
DRAM[55093] = 8'b11001001;
DRAM[55094] = 8'b11000111;
DRAM[55095] = 8'b11000101;
DRAM[55096] = 8'b10111111;
DRAM[55097] = 8'b11000111;
DRAM[55098] = 8'b11001001;
DRAM[55099] = 8'b11000101;
DRAM[55100] = 8'b11000110;
DRAM[55101] = 8'b11001001;
DRAM[55102] = 8'b11000000;
DRAM[55103] = 8'b10110001;
DRAM[55104] = 8'b10011110;
DRAM[55105] = 8'b10011100;
DRAM[55106] = 8'b10011101;
DRAM[55107] = 8'b10100000;
DRAM[55108] = 8'b10100011;
DRAM[55109] = 8'b10100100;
DRAM[55110] = 8'b10100100;
DRAM[55111] = 8'b10100101;
DRAM[55112] = 8'b10010111;
DRAM[55113] = 8'b10100010;
DRAM[55114] = 8'b10101100;
DRAM[55115] = 8'b10101001;
DRAM[55116] = 8'b10011101;
DRAM[55117] = 8'b10010101;
DRAM[55118] = 8'b10010110;
DRAM[55119] = 8'b10011011;
DRAM[55120] = 8'b10010110;
DRAM[55121] = 8'b10001100;
DRAM[55122] = 8'b10010010;
DRAM[55123] = 8'b10011110;
DRAM[55124] = 8'b10100000;
DRAM[55125] = 8'b10100010;
DRAM[55126] = 8'b10100010;
DRAM[55127] = 8'b10011010;
DRAM[55128] = 8'b10010001;
DRAM[55129] = 8'b10011010;
DRAM[55130] = 8'b10010110;
DRAM[55131] = 8'b10001011;
DRAM[55132] = 8'b10000101;
DRAM[55133] = 8'b10000000;
DRAM[55134] = 8'b10000010;
DRAM[55135] = 8'b10001111;
DRAM[55136] = 8'b10000011;
DRAM[55137] = 8'b1110011;
DRAM[55138] = 8'b1110101;
DRAM[55139] = 8'b1110000;
DRAM[55140] = 8'b1110100;
DRAM[55141] = 8'b1111100;
DRAM[55142] = 8'b1110110;
DRAM[55143] = 8'b1111111;
DRAM[55144] = 8'b10000000;
DRAM[55145] = 8'b1100100;
DRAM[55146] = 8'b1101011;
DRAM[55147] = 8'b1110111;
DRAM[55148] = 8'b1100101;
DRAM[55149] = 8'b1011110;
DRAM[55150] = 8'b1011101;
DRAM[55151] = 8'b1001001;
DRAM[55152] = 8'b1100010;
DRAM[55153] = 8'b1011010;
DRAM[55154] = 8'b1011001;
DRAM[55155] = 8'b1100001;
DRAM[55156] = 8'b1010101;
DRAM[55157] = 8'b1011100;
DRAM[55158] = 8'b1000000;
DRAM[55159] = 8'b1011110;
DRAM[55160] = 8'b1110000;
DRAM[55161] = 8'b1100110;
DRAM[55162] = 8'b1100001;
DRAM[55163] = 8'b1100011;
DRAM[55164] = 8'b1100101;
DRAM[55165] = 8'b1100010;
DRAM[55166] = 8'b1100000;
DRAM[55167] = 8'b1100010;
DRAM[55168] = 8'b1010100;
DRAM[55169] = 8'b1010011;
DRAM[55170] = 8'b1011100;
DRAM[55171] = 8'b1100000;
DRAM[55172] = 8'b1011111;
DRAM[55173] = 8'b1100101;
DRAM[55174] = 8'b1101001;
DRAM[55175] = 8'b1011111;
DRAM[55176] = 8'b1101000;
DRAM[55177] = 8'b1100011;
DRAM[55178] = 8'b1011110;
DRAM[55179] = 8'b1010011;
DRAM[55180] = 8'b1010000;
DRAM[55181] = 8'b1100010;
DRAM[55182] = 8'b1110001;
DRAM[55183] = 8'b1101011;
DRAM[55184] = 8'b1100000;
DRAM[55185] = 8'b1011000;
DRAM[55186] = 8'b1011000;
DRAM[55187] = 8'b1100111;
DRAM[55188] = 8'b1110011;
DRAM[55189] = 8'b1110001;
DRAM[55190] = 8'b1101000;
DRAM[55191] = 8'b1100010;
DRAM[55192] = 8'b1101100;
DRAM[55193] = 8'b1110111;
DRAM[55194] = 8'b1110111;
DRAM[55195] = 8'b10001000;
DRAM[55196] = 8'b1111011;
DRAM[55197] = 8'b10000111;
DRAM[55198] = 8'b10000010;
DRAM[55199] = 8'b10001101;
DRAM[55200] = 8'b10001010;
DRAM[55201] = 8'b10001100;
DRAM[55202] = 8'b10001111;
DRAM[55203] = 8'b10010000;
DRAM[55204] = 8'b10001111;
DRAM[55205] = 8'b10001110;
DRAM[55206] = 8'b10001110;
DRAM[55207] = 8'b10001111;
DRAM[55208] = 8'b10010010;
DRAM[55209] = 8'b10011000;
DRAM[55210] = 8'b10010101;
DRAM[55211] = 8'b10010101;
DRAM[55212] = 8'b10011111;
DRAM[55213] = 8'b10100001;
DRAM[55214] = 8'b10100001;
DRAM[55215] = 8'b10101001;
DRAM[55216] = 8'b10100011;
DRAM[55217] = 8'b10101001;
DRAM[55218] = 8'b10110010;
DRAM[55219] = 8'b10111010;
DRAM[55220] = 8'b11000001;
DRAM[55221] = 8'b11001001;
DRAM[55222] = 8'b11010010;
DRAM[55223] = 8'b11011000;
DRAM[55224] = 8'b11010110;
DRAM[55225] = 8'b11011110;
DRAM[55226] = 8'b11100100;
DRAM[55227] = 8'b11100100;
DRAM[55228] = 8'b11100010;
DRAM[55229] = 8'b11100101;
DRAM[55230] = 8'b11110001;
DRAM[55231] = 8'b11111101;
DRAM[55232] = 8'b11100101;
DRAM[55233] = 8'b11011101;
DRAM[55234] = 8'b11011001;
DRAM[55235] = 8'b11011011;
DRAM[55236] = 8'b11010101;
DRAM[55237] = 8'b11000011;
DRAM[55238] = 8'b10110010;
DRAM[55239] = 8'b10101001;
DRAM[55240] = 8'b10010011;
DRAM[55241] = 8'b10010100;
DRAM[55242] = 8'b10010100;
DRAM[55243] = 8'b10010001;
DRAM[55244] = 8'b10001010;
DRAM[55245] = 8'b10000100;
DRAM[55246] = 8'b10000001;
DRAM[55247] = 8'b10000000;
DRAM[55248] = 8'b1111010;
DRAM[55249] = 8'b1111101;
DRAM[55250] = 8'b1111100;
DRAM[55251] = 8'b1111000;
DRAM[55252] = 8'b1111000;
DRAM[55253] = 8'b1111011;
DRAM[55254] = 8'b1111011;
DRAM[55255] = 8'b1111000;
DRAM[55256] = 8'b1110111;
DRAM[55257] = 8'b1110110;
DRAM[55258] = 8'b1110011;
DRAM[55259] = 8'b1110001;
DRAM[55260] = 8'b1110000;
DRAM[55261] = 8'b1101111;
DRAM[55262] = 8'b1110000;
DRAM[55263] = 8'b1110000;
DRAM[55264] = 8'b1101110;
DRAM[55265] = 8'b1101110;
DRAM[55266] = 8'b1101110;
DRAM[55267] = 8'b1101111;
DRAM[55268] = 8'b1110000;
DRAM[55269] = 8'b1110001;
DRAM[55270] = 8'b1110010;
DRAM[55271] = 8'b1110011;
DRAM[55272] = 8'b1110001;
DRAM[55273] = 8'b1110001;
DRAM[55274] = 8'b1110001;
DRAM[55275] = 8'b1110001;
DRAM[55276] = 8'b1110000;
DRAM[55277] = 8'b1101111;
DRAM[55278] = 8'b1101110;
DRAM[55279] = 8'b1101101;
DRAM[55280] = 8'b1101101;
DRAM[55281] = 8'b1101101;
DRAM[55282] = 8'b1101101;
DRAM[55283] = 8'b1101101;
DRAM[55284] = 8'b1101100;
DRAM[55285] = 8'b1101011;
DRAM[55286] = 8'b1101010;
DRAM[55287] = 8'b1101001;
DRAM[55288] = 8'b1101001;
DRAM[55289] = 8'b1101001;
DRAM[55290] = 8'b1101010;
DRAM[55291] = 8'b1101010;
DRAM[55292] = 8'b1101011;
DRAM[55293] = 8'b1101100;
DRAM[55294] = 8'b1101101;
DRAM[55295] = 8'b1101101;
DRAM[55296] = 8'b10010100;
DRAM[55297] = 8'b10010101;
DRAM[55298] = 8'b10010110;
DRAM[55299] = 8'b10010111;
DRAM[55300] = 8'b10011001;
DRAM[55301] = 8'b10011011;
DRAM[55302] = 8'b10011100;
DRAM[55303] = 8'b10011100;
DRAM[55304] = 8'b10011101;
DRAM[55305] = 8'b10011110;
DRAM[55306] = 8'b10011111;
DRAM[55307] = 8'b10011111;
DRAM[55308] = 8'b10011101;
DRAM[55309] = 8'b10011101;
DRAM[55310] = 8'b10011110;
DRAM[55311] = 8'b10011111;
DRAM[55312] = 8'b10100000;
DRAM[55313] = 8'b10100110;
DRAM[55314] = 8'b10110101;
DRAM[55315] = 8'b11001010;
DRAM[55316] = 8'b11100000;
DRAM[55317] = 8'b11110010;
DRAM[55318] = 8'b11111101;
DRAM[55319] = 8'b11111111;
DRAM[55320] = 8'b11111011;
DRAM[55321] = 8'b11111100;
DRAM[55322] = 8'b11111100;
DRAM[55323] = 8'b11111100;
DRAM[55324] = 8'b11111100;
DRAM[55325] = 8'b11111011;
DRAM[55326] = 8'b11111010;
DRAM[55327] = 8'b11111001;
DRAM[55328] = 8'b11110110;
DRAM[55329] = 8'b11110101;
DRAM[55330] = 8'b11110100;
DRAM[55331] = 8'b11110010;
DRAM[55332] = 8'b11101111;
DRAM[55333] = 8'b11101110;
DRAM[55334] = 8'b11101101;
DRAM[55335] = 8'b11101101;
DRAM[55336] = 8'b11101101;
DRAM[55337] = 8'b11100111;
DRAM[55338] = 8'b11100010;
DRAM[55339] = 8'b11100011;
DRAM[55340] = 8'b11100111;
DRAM[55341] = 8'b11100111;
DRAM[55342] = 8'b11100000;
DRAM[55343] = 8'b11011001;
DRAM[55344] = 8'b11001110;
DRAM[55345] = 8'b11000111;
DRAM[55346] = 8'b10111111;
DRAM[55347] = 8'b10111100;
DRAM[55348] = 8'b11000001;
DRAM[55349] = 8'b11001010;
DRAM[55350] = 8'b11010100;
DRAM[55351] = 8'b11011010;
DRAM[55352] = 8'b11011000;
DRAM[55353] = 8'b11010101;
DRAM[55354] = 8'b11001111;
DRAM[55355] = 8'b11001011;
DRAM[55356] = 8'b11000110;
DRAM[55357] = 8'b11000001;
DRAM[55358] = 8'b10111011;
DRAM[55359] = 8'b10110111;
DRAM[55360] = 8'b10110110;
DRAM[55361] = 8'b10110000;
DRAM[55362] = 8'b10110011;
DRAM[55363] = 8'b10100110;
DRAM[55364] = 8'b10100100;
DRAM[55365] = 8'b10101010;
DRAM[55366] = 8'b10011101;
DRAM[55367] = 8'b10011101;
DRAM[55368] = 8'b10100111;
DRAM[55369] = 8'b10011011;
DRAM[55370] = 8'b10100000;
DRAM[55371] = 8'b10100010;
DRAM[55372] = 8'b10011000;
DRAM[55373] = 8'b10011101;
DRAM[55374] = 8'b10100000;
DRAM[55375] = 8'b10010001;
DRAM[55376] = 8'b10010010;
DRAM[55377] = 8'b10100000;
DRAM[55378] = 8'b10011110;
DRAM[55379] = 8'b10011000;
DRAM[55380] = 8'b10100010;
DRAM[55381] = 8'b10101000;
DRAM[55382] = 8'b10100000;
DRAM[55383] = 8'b10011000;
DRAM[55384] = 8'b10011100;
DRAM[55385] = 8'b10011111;
DRAM[55386] = 8'b10001110;
DRAM[55387] = 8'b10010010;
DRAM[55388] = 8'b10000010;
DRAM[55389] = 8'b10001111;
DRAM[55390] = 8'b10000011;
DRAM[55391] = 8'b10000100;
DRAM[55392] = 8'b10001111;
DRAM[55393] = 8'b1101110;
DRAM[55394] = 8'b1101101;
DRAM[55395] = 8'b1111110;
DRAM[55396] = 8'b1111100;
DRAM[55397] = 8'b1111010;
DRAM[55398] = 8'b10000000;
DRAM[55399] = 8'b1111011;
DRAM[55400] = 8'b1110110;
DRAM[55401] = 8'b1110000;
DRAM[55402] = 8'b1101111;
DRAM[55403] = 8'b1101111;
DRAM[55404] = 8'b1100101;
DRAM[55405] = 8'b1010110;
DRAM[55406] = 8'b1010101;
DRAM[55407] = 8'b1011110;
DRAM[55408] = 8'b1100010;
DRAM[55409] = 8'b1010100;
DRAM[55410] = 8'b1001111;
DRAM[55411] = 8'b1010110;
DRAM[55412] = 8'b1011001;
DRAM[55413] = 8'b1010000;
DRAM[55414] = 8'b1001001;
DRAM[55415] = 8'b1001001;
DRAM[55416] = 8'b1011110;
DRAM[55417] = 8'b1100100;
DRAM[55418] = 8'b1110100;
DRAM[55419] = 8'b1100001;
DRAM[55420] = 8'b1100000;
DRAM[55421] = 8'b1101010;
DRAM[55422] = 8'b1011011;
DRAM[55423] = 8'b1101100;
DRAM[55424] = 8'b1011010;
DRAM[55425] = 8'b1011000;
DRAM[55426] = 8'b1100001;
DRAM[55427] = 8'b1011000;
DRAM[55428] = 8'b1011010;
DRAM[55429] = 8'b1100101;
DRAM[55430] = 8'b1011011;
DRAM[55431] = 8'b1011010;
DRAM[55432] = 8'b1011100;
DRAM[55433] = 8'b1010101;
DRAM[55434] = 8'b1010010;
DRAM[55435] = 8'b1010111;
DRAM[55436] = 8'b1011101;
DRAM[55437] = 8'b1011101;
DRAM[55438] = 8'b1011100;
DRAM[55439] = 8'b1011100;
DRAM[55440] = 8'b1011010;
DRAM[55441] = 8'b1100110;
DRAM[55442] = 8'b1100110;
DRAM[55443] = 8'b1011000;
DRAM[55444] = 8'b1010101;
DRAM[55445] = 8'b1100011;
DRAM[55446] = 8'b1101011;
DRAM[55447] = 8'b1101001;
DRAM[55448] = 8'b1101001;
DRAM[55449] = 8'b1101101;
DRAM[55450] = 8'b1110110;
DRAM[55451] = 8'b1111111;
DRAM[55452] = 8'b1111111;
DRAM[55453] = 8'b1111100;
DRAM[55454] = 8'b10000001;
DRAM[55455] = 8'b10001010;
DRAM[55456] = 8'b10001101;
DRAM[55457] = 8'b10010000;
DRAM[55458] = 8'b10010010;
DRAM[55459] = 8'b10010001;
DRAM[55460] = 8'b10010001;
DRAM[55461] = 8'b10010010;
DRAM[55462] = 8'b10010111;
DRAM[55463] = 8'b10011011;
DRAM[55464] = 8'b10010001;
DRAM[55465] = 8'b10001111;
DRAM[55466] = 8'b10010000;
DRAM[55467] = 8'b10011000;
DRAM[55468] = 8'b10100011;
DRAM[55469] = 8'b10101010;
DRAM[55470] = 8'b10101000;
DRAM[55471] = 8'b10100101;
DRAM[55472] = 8'b10101011;
DRAM[55473] = 8'b10101101;
DRAM[55474] = 8'b10110000;
DRAM[55475] = 8'b10110011;
DRAM[55476] = 8'b10111000;
DRAM[55477] = 8'b11000010;
DRAM[55478] = 8'b11001110;
DRAM[55479] = 8'b11010111;
DRAM[55480] = 8'b11011011;
DRAM[55481] = 8'b11011001;
DRAM[55482] = 8'b11011000;
DRAM[55483] = 8'b11011101;
DRAM[55484] = 8'b11100110;
DRAM[55485] = 8'b11101110;
DRAM[55486] = 8'b11110001;
DRAM[55487] = 8'b11110001;
DRAM[55488] = 8'b11110011;
DRAM[55489] = 8'b11011011;
DRAM[55490] = 8'b11000010;
DRAM[55491] = 8'b10111001;
DRAM[55492] = 8'b10111000;
DRAM[55493] = 8'b10111000;
DRAM[55494] = 8'b10111010;
DRAM[55495] = 8'b10111101;
DRAM[55496] = 8'b10100000;
DRAM[55497] = 8'b10011011;
DRAM[55498] = 8'b10010100;
DRAM[55499] = 8'b10001101;
DRAM[55500] = 8'b10001000;
DRAM[55501] = 8'b10000101;
DRAM[55502] = 8'b10000101;
DRAM[55503] = 8'b10000101;
DRAM[55504] = 8'b1111110;
DRAM[55505] = 8'b1111101;
DRAM[55506] = 8'b1111100;
DRAM[55507] = 8'b1111011;
DRAM[55508] = 8'b1111010;
DRAM[55509] = 8'b1111001;
DRAM[55510] = 8'b1111001;
DRAM[55511] = 8'b1111001;
DRAM[55512] = 8'b1110111;
DRAM[55513] = 8'b1110101;
DRAM[55514] = 8'b1110011;
DRAM[55515] = 8'b1110010;
DRAM[55516] = 8'b1110010;
DRAM[55517] = 8'b1110001;
DRAM[55518] = 8'b1101111;
DRAM[55519] = 8'b1101101;
DRAM[55520] = 8'b1101101;
DRAM[55521] = 8'b1101101;
DRAM[55522] = 8'b1101101;
DRAM[55523] = 8'b1101101;
DRAM[55524] = 8'b1101110;
DRAM[55525] = 8'b1101111;
DRAM[55526] = 8'b1110000;
DRAM[55527] = 8'b1110000;
DRAM[55528] = 8'b1110000;
DRAM[55529] = 8'b1101111;
DRAM[55530] = 8'b1101110;
DRAM[55531] = 8'b1101110;
DRAM[55532] = 8'b1101101;
DRAM[55533] = 8'b1101101;
DRAM[55534] = 8'b1101110;
DRAM[55535] = 8'b1101110;
DRAM[55536] = 8'b1101100;
DRAM[55537] = 8'b1101100;
DRAM[55538] = 8'b1101011;
DRAM[55539] = 8'b1101010;
DRAM[55540] = 8'b1101010;
DRAM[55541] = 8'b1101001;
DRAM[55542] = 8'b1101000;
DRAM[55543] = 8'b1101000;
DRAM[55544] = 8'b1101000;
DRAM[55545] = 8'b1101000;
DRAM[55546] = 8'b1101001;
DRAM[55547] = 8'b1101010;
DRAM[55548] = 8'b1101010;
DRAM[55549] = 8'b1101011;
DRAM[55550] = 8'b1101100;
DRAM[55551] = 8'b1101100;
DRAM[55552] = 8'b10010011;
DRAM[55553] = 8'b10010100;
DRAM[55554] = 8'b10010101;
DRAM[55555] = 8'b10010111;
DRAM[55556] = 8'b10011000;
DRAM[55557] = 8'b10011010;
DRAM[55558] = 8'b10011011;
DRAM[55559] = 8'b10011100;
DRAM[55560] = 8'b10011101;
DRAM[55561] = 8'b10011110;
DRAM[55562] = 8'b10011111;
DRAM[55563] = 8'b10011111;
DRAM[55564] = 8'b10011110;
DRAM[55565] = 8'b10011101;
DRAM[55566] = 8'b10011111;
DRAM[55567] = 8'b10100000;
DRAM[55568] = 8'b10100001;
DRAM[55569] = 8'b10101000;
DRAM[55570] = 8'b10110111;
DRAM[55571] = 8'b11001101;
DRAM[55572] = 8'b11100100;
DRAM[55573] = 8'b11110101;
DRAM[55574] = 8'b11111100;
DRAM[55575] = 8'b11111110;
DRAM[55576] = 8'b11111100;
DRAM[55577] = 8'b11111100;
DRAM[55578] = 8'b11111101;
DRAM[55579] = 8'b11111100;
DRAM[55580] = 8'b11111100;
DRAM[55581] = 8'b11111011;
DRAM[55582] = 8'b11111001;
DRAM[55583] = 8'b11111001;
DRAM[55584] = 8'b11110011;
DRAM[55585] = 8'b11110001;
DRAM[55586] = 8'b11110000;
DRAM[55587] = 8'b11110000;
DRAM[55588] = 8'b11110010;
DRAM[55589] = 8'b11110100;
DRAM[55590] = 8'b11110101;
DRAM[55591] = 8'b11110110;
DRAM[55592] = 8'b11111000;
DRAM[55593] = 8'b11110000;
DRAM[55594] = 8'b11100111;
DRAM[55595] = 8'b11100010;
DRAM[55596] = 8'b11100001;
DRAM[55597] = 8'b11100000;
DRAM[55598] = 8'b11011011;
DRAM[55599] = 8'b11010110;
DRAM[55600] = 8'b11010111;
DRAM[55601] = 8'b11010011;
DRAM[55602] = 8'b11001111;
DRAM[55603] = 8'b11001100;
DRAM[55604] = 8'b11001101;
DRAM[55605] = 8'b11001110;
DRAM[55606] = 8'b11001111;
DRAM[55607] = 8'b11001111;
DRAM[55608] = 8'b11010110;
DRAM[55609] = 8'b11010010;
DRAM[55610] = 8'b11001100;
DRAM[55611] = 8'b11001000;
DRAM[55612] = 8'b11000110;
DRAM[55613] = 8'b11000101;
DRAM[55614] = 8'b11000011;
DRAM[55615] = 8'b11000001;
DRAM[55616] = 8'b11001000;
DRAM[55617] = 8'b10110011;
DRAM[55618] = 8'b10101110;
DRAM[55619] = 8'b10100001;
DRAM[55620] = 8'b10011100;
DRAM[55621] = 8'b10011110;
DRAM[55622] = 8'b10011010;
DRAM[55623] = 8'b10101010;
DRAM[55624] = 8'b10100011;
DRAM[55625] = 8'b10011100;
DRAM[55626] = 8'b10011011;
DRAM[55627] = 8'b10011010;
DRAM[55628] = 8'b10010101;
DRAM[55629] = 8'b10011010;
DRAM[55630] = 8'b10011111;
DRAM[55631] = 8'b10011010;
DRAM[55632] = 8'b10100100;
DRAM[55633] = 8'b10100100;
DRAM[55634] = 8'b10100010;
DRAM[55635] = 8'b10100111;
DRAM[55636] = 8'b10101000;
DRAM[55637] = 8'b10011000;
DRAM[55638] = 8'b10010000;
DRAM[55639] = 8'b10011100;
DRAM[55640] = 8'b10010110;
DRAM[55641] = 8'b10011010;
DRAM[55642] = 8'b10001101;
DRAM[55643] = 8'b10010000;
DRAM[55644] = 8'b10000001;
DRAM[55645] = 8'b10001011;
DRAM[55646] = 8'b1111110;
DRAM[55647] = 8'b1111100;
DRAM[55648] = 8'b10000110;
DRAM[55649] = 8'b1101010;
DRAM[55650] = 8'b1101001;
DRAM[55651] = 8'b1111001;
DRAM[55652] = 8'b1110111;
DRAM[55653] = 8'b1110101;
DRAM[55654] = 8'b1111100;
DRAM[55655] = 8'b1111001;
DRAM[55656] = 8'b1110001;
DRAM[55657] = 8'b1101100;
DRAM[55658] = 8'b1101011;
DRAM[55659] = 8'b1101011;
DRAM[55660] = 8'b1100010;
DRAM[55661] = 8'b1010101;
DRAM[55662] = 8'b1010100;
DRAM[55663] = 8'b1011100;
DRAM[55664] = 8'b1011111;
DRAM[55665] = 8'b1010101;
DRAM[55666] = 8'b1010011;
DRAM[55667] = 8'b1011010;
DRAM[55668] = 8'b1011011;
DRAM[55669] = 8'b1010010;
DRAM[55670] = 8'b1001100;
DRAM[55671] = 8'b1001110;
DRAM[55672] = 8'b1011101;
DRAM[55673] = 8'b1100101;
DRAM[55674] = 8'b1101010;
DRAM[55675] = 8'b1100000;
DRAM[55676] = 8'b1100100;
DRAM[55677] = 8'b1101010;
DRAM[55678] = 8'b1100000;
DRAM[55679] = 8'b1101000;
DRAM[55680] = 8'b1011010;
DRAM[55681] = 8'b1010111;
DRAM[55682] = 8'b1100000;
DRAM[55683] = 8'b1011000;
DRAM[55684] = 8'b1011001;
DRAM[55685] = 8'b1100010;
DRAM[55686] = 8'b1010111;
DRAM[55687] = 8'b1010111;
DRAM[55688] = 8'b1010101;
DRAM[55689] = 8'b1010000;
DRAM[55690] = 8'b1001111;
DRAM[55691] = 8'b1010100;
DRAM[55692] = 8'b1010111;
DRAM[55693] = 8'b1011000;
DRAM[55694] = 8'b1011011;
DRAM[55695] = 8'b1011111;
DRAM[55696] = 8'b1011001;
DRAM[55697] = 8'b1011101;
DRAM[55698] = 8'b1011111;
DRAM[55699] = 8'b1011111;
DRAM[55700] = 8'b1011111;
DRAM[55701] = 8'b1100011;
DRAM[55702] = 8'b1101001;
DRAM[55703] = 8'b1101101;
DRAM[55704] = 8'b1101110;
DRAM[55705] = 8'b1110001;
DRAM[55706] = 8'b1111001;
DRAM[55707] = 8'b10000001;
DRAM[55708] = 8'b10000001;
DRAM[55709] = 8'b1111011;
DRAM[55710] = 8'b1111011;
DRAM[55711] = 8'b10000000;
DRAM[55712] = 8'b10000101;
DRAM[55713] = 8'b10001001;
DRAM[55714] = 8'b10001110;
DRAM[55715] = 8'b10010001;
DRAM[55716] = 8'b10010010;
DRAM[55717] = 8'b10010011;
DRAM[55718] = 8'b10010101;
DRAM[55719] = 8'b10010111;
DRAM[55720] = 8'b10011000;
DRAM[55721] = 8'b10011100;
DRAM[55722] = 8'b10011110;
DRAM[55723] = 8'b10011100;
DRAM[55724] = 8'b10011010;
DRAM[55725] = 8'b10011101;
DRAM[55726] = 8'b10100111;
DRAM[55727] = 8'b10110000;
DRAM[55728] = 8'b10101111;
DRAM[55729] = 8'b10110000;
DRAM[55730] = 8'b10110010;
DRAM[55731] = 8'b10110011;
DRAM[55732] = 8'b10110101;
DRAM[55733] = 8'b10111011;
DRAM[55734] = 8'b11000011;
DRAM[55735] = 8'b11001001;
DRAM[55736] = 8'b11011000;
DRAM[55737] = 8'b11011100;
DRAM[55738] = 8'b11100001;
DRAM[55739] = 8'b11100111;
DRAM[55740] = 8'b11101011;
DRAM[55741] = 8'b11101110;
DRAM[55742] = 8'b11110001;
DRAM[55743] = 8'b11110011;
DRAM[55744] = 8'b11100110;
DRAM[55745] = 8'b11010100;
DRAM[55746] = 8'b10111101;
DRAM[55747] = 8'b10101100;
DRAM[55748] = 8'b10011110;
DRAM[55749] = 8'b10010011;
DRAM[55750] = 8'b10001111;
DRAM[55751] = 8'b10010010;
DRAM[55752] = 8'b10010100;
DRAM[55753] = 8'b10010011;
DRAM[55754] = 8'b10010000;
DRAM[55755] = 8'b10001101;
DRAM[55756] = 8'b10001001;
DRAM[55757] = 8'b10000110;
DRAM[55758] = 8'b10000100;
DRAM[55759] = 8'b10000011;
DRAM[55760] = 8'b1111011;
DRAM[55761] = 8'b1111010;
DRAM[55762] = 8'b1111010;
DRAM[55763] = 8'b1111001;
DRAM[55764] = 8'b1111001;
DRAM[55765] = 8'b1111001;
DRAM[55766] = 8'b1111010;
DRAM[55767] = 8'b1111010;
DRAM[55768] = 8'b1111001;
DRAM[55769] = 8'b1110111;
DRAM[55770] = 8'b1110100;
DRAM[55771] = 8'b1110011;
DRAM[55772] = 8'b1110011;
DRAM[55773] = 8'b1110010;
DRAM[55774] = 8'b1110000;
DRAM[55775] = 8'b1101110;
DRAM[55776] = 8'b1101110;
DRAM[55777] = 8'b1101110;
DRAM[55778] = 8'b1101101;
DRAM[55779] = 8'b1101101;
DRAM[55780] = 8'b1101101;
DRAM[55781] = 8'b1101110;
DRAM[55782] = 8'b1101111;
DRAM[55783] = 8'b1101111;
DRAM[55784] = 8'b1101111;
DRAM[55785] = 8'b1101110;
DRAM[55786] = 8'b1101110;
DRAM[55787] = 8'b1101101;
DRAM[55788] = 8'b1101100;
DRAM[55789] = 8'b1101100;
DRAM[55790] = 8'b1101101;
DRAM[55791] = 8'b1101101;
DRAM[55792] = 8'b1101100;
DRAM[55793] = 8'b1101100;
DRAM[55794] = 8'b1101011;
DRAM[55795] = 8'b1101010;
DRAM[55796] = 8'b1101010;
DRAM[55797] = 8'b1101001;
DRAM[55798] = 8'b1101000;
DRAM[55799] = 8'b1101000;
DRAM[55800] = 8'b1101000;
DRAM[55801] = 8'b1101000;
DRAM[55802] = 8'b1101001;
DRAM[55803] = 8'b1101010;
DRAM[55804] = 8'b1101010;
DRAM[55805] = 8'b1101011;
DRAM[55806] = 8'b1101100;
DRAM[55807] = 8'b1101100;
DRAM[55808] = 8'b10010010;
DRAM[55809] = 8'b10010011;
DRAM[55810] = 8'b10010100;
DRAM[55811] = 8'b10010110;
DRAM[55812] = 8'b10010111;
DRAM[55813] = 8'b10011001;
DRAM[55814] = 8'b10011010;
DRAM[55815] = 8'b10011011;
DRAM[55816] = 8'b10011100;
DRAM[55817] = 8'b10011110;
DRAM[55818] = 8'b10100000;
DRAM[55819] = 8'b10100000;
DRAM[55820] = 8'b10011111;
DRAM[55821] = 8'b10011111;
DRAM[55822] = 8'b10100000;
DRAM[55823] = 8'b10100010;
DRAM[55824] = 8'b10100100;
DRAM[55825] = 8'b10101100;
DRAM[55826] = 8'b10111100;
DRAM[55827] = 8'b11010011;
DRAM[55828] = 8'b11101010;
DRAM[55829] = 8'b11111000;
DRAM[55830] = 8'b11111100;
DRAM[55831] = 8'b11111011;
DRAM[55832] = 8'b11111101;
DRAM[55833] = 8'b11111101;
DRAM[55834] = 8'b11111101;
DRAM[55835] = 8'b11111101;
DRAM[55836] = 8'b11111100;
DRAM[55837] = 8'b11111010;
DRAM[55838] = 8'b11111001;
DRAM[55839] = 8'b11111000;
DRAM[55840] = 8'b11110110;
DRAM[55841] = 8'b11110011;
DRAM[55842] = 8'b11101111;
DRAM[55843] = 8'b11110000;
DRAM[55844] = 8'b11110011;
DRAM[55845] = 8'b11110110;
DRAM[55846] = 8'b11110110;
DRAM[55847] = 8'b11110101;
DRAM[55848] = 8'b11100111;
DRAM[55849] = 8'b11100100;
DRAM[55850] = 8'b11100001;
DRAM[55851] = 8'b11011111;
DRAM[55852] = 8'b11011111;
DRAM[55853] = 8'b11011110;
DRAM[55854] = 8'b11011011;
DRAM[55855] = 8'b11011001;
DRAM[55856] = 8'b11010011;
DRAM[55857] = 8'b11010100;
DRAM[55858] = 8'b11010110;
DRAM[55859] = 8'b11011001;
DRAM[55860] = 8'b11011010;
DRAM[55861] = 8'b11011000;
DRAM[55862] = 8'b11010010;
DRAM[55863] = 8'b11001110;
DRAM[55864] = 8'b11001101;
DRAM[55865] = 8'b11001000;
DRAM[55866] = 8'b11000011;
DRAM[55867] = 8'b11000000;
DRAM[55868] = 8'b11000001;
DRAM[55869] = 8'b11000011;
DRAM[55870] = 8'b11000101;
DRAM[55871] = 8'b11000101;
DRAM[55872] = 8'b10111110;
DRAM[55873] = 8'b10101111;
DRAM[55874] = 8'b10111010;
DRAM[55875] = 8'b10111101;
DRAM[55876] = 8'b10110111;
DRAM[55877] = 8'b10101000;
DRAM[55878] = 8'b10010111;
DRAM[55879] = 8'b10100100;
DRAM[55880] = 8'b10011011;
DRAM[55881] = 8'b10011111;
DRAM[55882] = 8'b10011100;
DRAM[55883] = 8'b10011001;
DRAM[55884] = 8'b10011100;
DRAM[55885] = 8'b10011010;
DRAM[55886] = 8'b10011000;
DRAM[55887] = 8'b10011110;
DRAM[55888] = 8'b10011100;
DRAM[55889] = 8'b10011111;
DRAM[55890] = 8'b10100000;
DRAM[55891] = 8'b10100011;
DRAM[55892] = 8'b10100001;
DRAM[55893] = 8'b10001111;
DRAM[55894] = 8'b10001011;
DRAM[55895] = 8'b10011011;
DRAM[55896] = 8'b10010101;
DRAM[55897] = 8'b10011001;
DRAM[55898] = 8'b10010001;
DRAM[55899] = 8'b10010011;
DRAM[55900] = 8'b10001000;
DRAM[55901] = 8'b10001100;
DRAM[55902] = 8'b10000000;
DRAM[55903] = 8'b1111100;
DRAM[55904] = 8'b1111101;
DRAM[55905] = 8'b1101010;
DRAM[55906] = 8'b1101011;
DRAM[55907] = 8'b1110110;
DRAM[55908] = 8'b1110100;
DRAM[55909] = 8'b1110100;
DRAM[55910] = 8'b1111010;
DRAM[55911] = 8'b1111011;
DRAM[55912] = 8'b1101110;
DRAM[55913] = 8'b1101010;
DRAM[55914] = 8'b1101001;
DRAM[55915] = 8'b1101001;
DRAM[55916] = 8'b1100010;
DRAM[55917] = 8'b1010111;
DRAM[55918] = 8'b1010110;
DRAM[55919] = 8'b1011100;
DRAM[55920] = 8'b1011011;
DRAM[55921] = 8'b1010111;
DRAM[55922] = 8'b1011001;
DRAM[55923] = 8'b1011111;
DRAM[55924] = 8'b1011110;
DRAM[55925] = 8'b1010100;
DRAM[55926] = 8'b1010000;
DRAM[55927] = 8'b1010010;
DRAM[55928] = 8'b1011011;
DRAM[55929] = 8'b1101000;
DRAM[55930] = 8'b1011111;
DRAM[55931] = 8'b1100010;
DRAM[55932] = 8'b1101011;
DRAM[55933] = 8'b1101000;
DRAM[55934] = 8'b1101001;
DRAM[55935] = 8'b1100110;
DRAM[55936] = 8'b1011111;
DRAM[55937] = 8'b1011010;
DRAM[55938] = 8'b1100010;
DRAM[55939] = 8'b1011010;
DRAM[55940] = 8'b1011010;
DRAM[55941] = 8'b1100001;
DRAM[55942] = 8'b1010101;
DRAM[55943] = 8'b1010101;
DRAM[55944] = 8'b1010100;
DRAM[55945] = 8'b1010100;
DRAM[55946] = 8'b1010111;
DRAM[55947] = 8'b1011001;
DRAM[55948] = 8'b1010110;
DRAM[55949] = 8'b1010100;
DRAM[55950] = 8'b1011010;
DRAM[55951] = 8'b1100011;
DRAM[55952] = 8'b1011101;
DRAM[55953] = 8'b1011000;
DRAM[55954] = 8'b1011011;
DRAM[55955] = 8'b1100100;
DRAM[55956] = 8'b1100110;
DRAM[55957] = 8'b1100010;
DRAM[55958] = 8'b1100011;
DRAM[55959] = 8'b1101010;
DRAM[55960] = 8'b1110000;
DRAM[55961] = 8'b1110010;
DRAM[55962] = 8'b1111001;
DRAM[55963] = 8'b10000001;
DRAM[55964] = 8'b10000010;
DRAM[55965] = 8'b1111101;
DRAM[55966] = 8'b1111001;
DRAM[55967] = 8'b1111001;
DRAM[55968] = 8'b1111101;
DRAM[55969] = 8'b10000011;
DRAM[55970] = 8'b10001011;
DRAM[55971] = 8'b10010001;
DRAM[55972] = 8'b10010100;
DRAM[55973] = 8'b10010101;
DRAM[55974] = 8'b10010110;
DRAM[55975] = 8'b10010110;
DRAM[55976] = 8'b10100000;
DRAM[55977] = 8'b10100011;
DRAM[55978] = 8'b10100100;
DRAM[55979] = 8'b10100001;
DRAM[55980] = 8'b10011100;
DRAM[55981] = 8'b10011101;
DRAM[55982] = 8'b10100100;
DRAM[55983] = 8'b10101100;
DRAM[55984] = 8'b10101111;
DRAM[55985] = 8'b10110001;
DRAM[55986] = 8'b10110011;
DRAM[55987] = 8'b10110101;
DRAM[55988] = 8'b10110101;
DRAM[55989] = 8'b10110111;
DRAM[55990] = 8'b10111001;
DRAM[55991] = 8'b10111100;
DRAM[55992] = 8'b11001110;
DRAM[55993] = 8'b11010111;
DRAM[55994] = 8'b11100100;
DRAM[55995] = 8'b11101100;
DRAM[55996] = 8'b11101110;
DRAM[55997] = 8'b11110000;
DRAM[55998] = 8'b11110011;
DRAM[55999] = 8'b11110110;
DRAM[56000] = 8'b11101110;
DRAM[56001] = 8'b11000111;
DRAM[56002] = 8'b10011110;
DRAM[56003] = 8'b10010001;
DRAM[56004] = 8'b10011001;
DRAM[56005] = 8'b10011100;
DRAM[56006] = 8'b10001111;
DRAM[56007] = 8'b10000000;
DRAM[56008] = 8'b10001000;
DRAM[56009] = 8'b10001001;
DRAM[56010] = 8'b10001011;
DRAM[56011] = 8'b10001011;
DRAM[56012] = 8'b10001010;
DRAM[56013] = 8'b10000111;
DRAM[56014] = 8'b10000100;
DRAM[56015] = 8'b10000001;
DRAM[56016] = 8'b1111001;
DRAM[56017] = 8'b1111000;
DRAM[56018] = 8'b1111000;
DRAM[56019] = 8'b1111000;
DRAM[56020] = 8'b1111000;
DRAM[56021] = 8'b1111001;
DRAM[56022] = 8'b1111010;
DRAM[56023] = 8'b1111011;
DRAM[56024] = 8'b1111010;
DRAM[56025] = 8'b1110111;
DRAM[56026] = 8'b1110101;
DRAM[56027] = 8'b1110100;
DRAM[56028] = 8'b1110100;
DRAM[56029] = 8'b1110011;
DRAM[56030] = 8'b1110001;
DRAM[56031] = 8'b1101111;
DRAM[56032] = 8'b1101111;
DRAM[56033] = 8'b1101110;
DRAM[56034] = 8'b1101110;
DRAM[56035] = 8'b1101101;
DRAM[56036] = 8'b1101101;
DRAM[56037] = 8'b1101101;
DRAM[56038] = 8'b1101101;
DRAM[56039] = 8'b1101110;
DRAM[56040] = 8'b1101110;
DRAM[56041] = 8'b1101101;
DRAM[56042] = 8'b1101100;
DRAM[56043] = 8'b1101011;
DRAM[56044] = 8'b1101011;
DRAM[56045] = 8'b1101011;
DRAM[56046] = 8'b1101011;
DRAM[56047] = 8'b1101011;
DRAM[56048] = 8'b1101100;
DRAM[56049] = 8'b1101100;
DRAM[56050] = 8'b1101011;
DRAM[56051] = 8'b1101010;
DRAM[56052] = 8'b1101010;
DRAM[56053] = 8'b1101001;
DRAM[56054] = 8'b1101000;
DRAM[56055] = 8'b1101000;
DRAM[56056] = 8'b1101000;
DRAM[56057] = 8'b1101000;
DRAM[56058] = 8'b1101001;
DRAM[56059] = 8'b1101010;
DRAM[56060] = 8'b1101010;
DRAM[56061] = 8'b1101011;
DRAM[56062] = 8'b1101100;
DRAM[56063] = 8'b1101100;
DRAM[56064] = 8'b10010001;
DRAM[56065] = 8'b10010001;
DRAM[56066] = 8'b10010010;
DRAM[56067] = 8'b10010100;
DRAM[56068] = 8'b10010110;
DRAM[56069] = 8'b10010111;
DRAM[56070] = 8'b10011000;
DRAM[56071] = 8'b10011001;
DRAM[56072] = 8'b10011100;
DRAM[56073] = 8'b10011101;
DRAM[56074] = 8'b10011111;
DRAM[56075] = 8'b10100000;
DRAM[56076] = 8'b10011111;
DRAM[56077] = 8'b10011111;
DRAM[56078] = 8'b10100001;
DRAM[56079] = 8'b10100011;
DRAM[56080] = 8'b10101000;
DRAM[56081] = 8'b10110001;
DRAM[56082] = 8'b11000011;
DRAM[56083] = 8'b11011011;
DRAM[56084] = 8'b11110001;
DRAM[56085] = 8'b11111100;
DRAM[56086] = 8'b11111100;
DRAM[56087] = 8'b11111000;
DRAM[56088] = 8'b11111110;
DRAM[56089] = 8'b11111101;
DRAM[56090] = 8'b11111101;
DRAM[56091] = 8'b11111100;
DRAM[56092] = 8'b11111011;
DRAM[56093] = 8'b11111001;
DRAM[56094] = 8'b11110111;
DRAM[56095] = 8'b11110110;
DRAM[56096] = 8'b11111011;
DRAM[56097] = 8'b11110111;
DRAM[56098] = 8'b11110011;
DRAM[56099] = 8'b11110011;
DRAM[56100] = 8'b11110100;
DRAM[56101] = 8'b11110010;
DRAM[56102] = 8'b11101101;
DRAM[56103] = 8'b11101000;
DRAM[56104] = 8'b11011010;
DRAM[56105] = 8'b11011101;
DRAM[56106] = 8'b11100001;
DRAM[56107] = 8'b11100100;
DRAM[56108] = 8'b11100100;
DRAM[56109] = 8'b11100010;
DRAM[56110] = 8'b11011110;
DRAM[56111] = 8'b11011100;
DRAM[56112] = 8'b11010010;
DRAM[56113] = 8'b11010011;
DRAM[56114] = 8'b11010111;
DRAM[56115] = 8'b11011011;
DRAM[56116] = 8'b11011100;
DRAM[56117] = 8'b11011001;
DRAM[56118] = 8'b11010011;
DRAM[56119] = 8'b11001111;
DRAM[56120] = 8'b11000100;
DRAM[56121] = 8'b11000001;
DRAM[56122] = 8'b10111100;
DRAM[56123] = 8'b10111011;
DRAM[56124] = 8'b10111011;
DRAM[56125] = 8'b10111101;
DRAM[56126] = 8'b10111110;
DRAM[56127] = 8'b10111110;
DRAM[56128] = 8'b11000001;
DRAM[56129] = 8'b10110100;
DRAM[56130] = 8'b10111000;
DRAM[56131] = 8'b10110010;
DRAM[56132] = 8'b10101100;
DRAM[56133] = 8'b10101010;
DRAM[56134] = 8'b10100100;
DRAM[56135] = 8'b10110010;
DRAM[56136] = 8'b10010000;
DRAM[56137] = 8'b10011111;
DRAM[56138] = 8'b10011111;
DRAM[56139] = 8'b10100000;
DRAM[56140] = 8'b10101000;
DRAM[56141] = 8'b10011100;
DRAM[56142] = 8'b10010000;
DRAM[56143] = 8'b10011011;
DRAM[56144] = 8'b10001101;
DRAM[56145] = 8'b10100000;
DRAM[56146] = 8'b10100001;
DRAM[56147] = 8'b10010100;
DRAM[56148] = 8'b10010011;
DRAM[56149] = 8'b10010100;
DRAM[56150] = 8'b10001111;
DRAM[56151] = 8'b10001111;
DRAM[56152] = 8'b10010100;
DRAM[56153] = 8'b10010111;
DRAM[56154] = 8'b10010011;
DRAM[56155] = 8'b10010000;
DRAM[56156] = 8'b10001011;
DRAM[56157] = 8'b10001101;
DRAM[56158] = 8'b10000110;
DRAM[56159] = 8'b1111111;
DRAM[56160] = 8'b1111010;
DRAM[56161] = 8'b1110010;
DRAM[56162] = 8'b1110010;
DRAM[56163] = 8'b1111000;
DRAM[56164] = 8'b1111000;
DRAM[56165] = 8'b1111000;
DRAM[56166] = 8'b1111101;
DRAM[56167] = 8'b10000010;
DRAM[56168] = 8'b1101111;
DRAM[56169] = 8'b1101011;
DRAM[56170] = 8'b1101010;
DRAM[56171] = 8'b1101010;
DRAM[56172] = 8'b1100100;
DRAM[56173] = 8'b1011100;
DRAM[56174] = 8'b1011011;
DRAM[56175] = 8'b1011111;
DRAM[56176] = 8'b1011001;
DRAM[56177] = 8'b1011010;
DRAM[56178] = 8'b1011111;
DRAM[56179] = 8'b1100011;
DRAM[56180] = 8'b1011111;
DRAM[56181] = 8'b1010101;
DRAM[56182] = 8'b1010001;
DRAM[56183] = 8'b1010011;
DRAM[56184] = 8'b1010110;
DRAM[56185] = 8'b1101010;
DRAM[56186] = 8'b1011100;
DRAM[56187] = 8'b1100111;
DRAM[56188] = 8'b1101111;
DRAM[56189] = 8'b1100100;
DRAM[56190] = 8'b1110000;
DRAM[56191] = 8'b1101011;
DRAM[56192] = 8'b1100111;
DRAM[56193] = 8'b1100000;
DRAM[56194] = 8'b1100111;
DRAM[56195] = 8'b1011111;
DRAM[56196] = 8'b1011110;
DRAM[56197] = 8'b1100011;
DRAM[56198] = 8'b1010110;
DRAM[56199] = 8'b1011001;
DRAM[56200] = 8'b1010100;
DRAM[56201] = 8'b1011000;
DRAM[56202] = 8'b1011111;
DRAM[56203] = 8'b1011111;
DRAM[56204] = 8'b1010111;
DRAM[56205] = 8'b1010000;
DRAM[56206] = 8'b1010100;
DRAM[56207] = 8'b1011101;
DRAM[56208] = 8'b1100000;
DRAM[56209] = 8'b1011101;
DRAM[56210] = 8'b1011101;
DRAM[56211] = 8'b1100001;
DRAM[56212] = 8'b1100011;
DRAM[56213] = 8'b1100010;
DRAM[56214] = 8'b1100000;
DRAM[56215] = 8'b1100001;
DRAM[56216] = 8'b1101111;
DRAM[56217] = 8'b1110001;
DRAM[56218] = 8'b1110110;
DRAM[56219] = 8'b1111101;
DRAM[56220] = 8'b10000001;
DRAM[56221] = 8'b10000000;
DRAM[56222] = 8'b1111101;
DRAM[56223] = 8'b1111010;
DRAM[56224] = 8'b1111100;
DRAM[56225] = 8'b10000000;
DRAM[56226] = 8'b10000111;
DRAM[56227] = 8'b10001110;
DRAM[56228] = 8'b10010011;
DRAM[56229] = 8'b10010110;
DRAM[56230] = 8'b10011000;
DRAM[56231] = 8'b10011001;
DRAM[56232] = 8'b10100010;
DRAM[56233] = 8'b10011111;
DRAM[56234] = 8'b10011110;
DRAM[56235] = 8'b10100011;
DRAM[56236] = 8'b10101001;
DRAM[56237] = 8'b10101011;
DRAM[56238] = 8'b10100101;
DRAM[56239] = 8'b10011111;
DRAM[56240] = 8'b10101100;
DRAM[56241] = 8'b10101111;
DRAM[56242] = 8'b10110011;
DRAM[56243] = 8'b10110111;
DRAM[56244] = 8'b10111001;
DRAM[56245] = 8'b10111010;
DRAM[56246] = 8'b10111010;
DRAM[56247] = 8'b10111010;
DRAM[56248] = 8'b11000011;
DRAM[56249] = 8'b11001100;
DRAM[56250] = 8'b11011010;
DRAM[56251] = 8'b11100110;
DRAM[56252] = 8'b11101110;
DRAM[56253] = 8'b11110011;
DRAM[56254] = 8'b11110111;
DRAM[56255] = 8'b11111001;
DRAM[56256] = 8'b11110001;
DRAM[56257] = 8'b11100111;
DRAM[56258] = 8'b11010011;
DRAM[56259] = 8'b10111000;
DRAM[56260] = 8'b10011100;
DRAM[56261] = 8'b10001011;
DRAM[56262] = 8'b10001001;
DRAM[56263] = 8'b10001110;
DRAM[56264] = 8'b10000011;
DRAM[56265] = 8'b10000101;
DRAM[56266] = 8'b10000111;
DRAM[56267] = 8'b10001001;
DRAM[56268] = 8'b10001001;
DRAM[56269] = 8'b10000111;
DRAM[56270] = 8'b10000100;
DRAM[56271] = 8'b10000010;
DRAM[56272] = 8'b1111011;
DRAM[56273] = 8'b1111010;
DRAM[56274] = 8'b1111001;
DRAM[56275] = 8'b1111001;
DRAM[56276] = 8'b1111000;
DRAM[56277] = 8'b1111001;
DRAM[56278] = 8'b1111001;
DRAM[56279] = 8'b1111010;
DRAM[56280] = 8'b1111001;
DRAM[56281] = 8'b1110111;
DRAM[56282] = 8'b1110101;
DRAM[56283] = 8'b1110100;
DRAM[56284] = 8'b1110100;
DRAM[56285] = 8'b1110011;
DRAM[56286] = 8'b1110000;
DRAM[56287] = 8'b1101110;
DRAM[56288] = 8'b1110000;
DRAM[56289] = 8'b1101111;
DRAM[56290] = 8'b1101110;
DRAM[56291] = 8'b1101101;
DRAM[56292] = 8'b1101100;
DRAM[56293] = 8'b1101100;
DRAM[56294] = 8'b1101100;
DRAM[56295] = 8'b1101100;
DRAM[56296] = 8'b1101100;
DRAM[56297] = 8'b1101100;
DRAM[56298] = 8'b1101011;
DRAM[56299] = 8'b1101010;
DRAM[56300] = 8'b1101001;
DRAM[56301] = 8'b1101001;
DRAM[56302] = 8'b1101010;
DRAM[56303] = 8'b1101010;
DRAM[56304] = 8'b1101011;
DRAM[56305] = 8'b1101011;
DRAM[56306] = 8'b1101011;
DRAM[56307] = 8'b1101010;
DRAM[56308] = 8'b1101010;
DRAM[56309] = 8'b1101001;
DRAM[56310] = 8'b1101001;
DRAM[56311] = 8'b1101001;
DRAM[56312] = 8'b1101001;
DRAM[56313] = 8'b1101001;
DRAM[56314] = 8'b1101001;
DRAM[56315] = 8'b1101010;
DRAM[56316] = 8'b1101010;
DRAM[56317] = 8'b1101011;
DRAM[56318] = 8'b1101011;
DRAM[56319] = 8'b1101011;
DRAM[56320] = 8'b10001111;
DRAM[56321] = 8'b10010000;
DRAM[56322] = 8'b10010001;
DRAM[56323] = 8'b10010010;
DRAM[56324] = 8'b10010100;
DRAM[56325] = 8'b10010110;
DRAM[56326] = 8'b10010111;
DRAM[56327] = 8'b10010111;
DRAM[56328] = 8'b10011010;
DRAM[56329] = 8'b10011100;
DRAM[56330] = 8'b10011110;
DRAM[56331] = 8'b10011111;
DRAM[56332] = 8'b10011111;
DRAM[56333] = 8'b10100000;
DRAM[56334] = 8'b10100010;
DRAM[56335] = 8'b10100100;
DRAM[56336] = 8'b10101011;
DRAM[56337] = 8'b10110111;
DRAM[56338] = 8'b11001100;
DRAM[56339] = 8'b11100100;
DRAM[56340] = 8'b11110110;
DRAM[56341] = 8'b11111101;
DRAM[56342] = 8'b11111100;
DRAM[56343] = 8'b11111000;
DRAM[56344] = 8'b11111101;
DRAM[56345] = 8'b11111101;
DRAM[56346] = 8'b11111101;
DRAM[56347] = 8'b11111011;
DRAM[56348] = 8'b11111001;
DRAM[56349] = 8'b11110111;
DRAM[56350] = 8'b11110101;
DRAM[56351] = 8'b11110100;
DRAM[56352] = 8'b11110100;
DRAM[56353] = 8'b11110011;
DRAM[56354] = 8'b11110011;
DRAM[56355] = 8'b11110100;
DRAM[56356] = 8'b11110100;
DRAM[56357] = 8'b11110000;
DRAM[56358] = 8'b11101001;
DRAM[56359] = 8'b11100100;
DRAM[56360] = 8'b11101100;
DRAM[56361] = 8'b11101100;
DRAM[56362] = 8'b11101011;
DRAM[56363] = 8'b11101010;
DRAM[56364] = 8'b11100111;
DRAM[56365] = 8'b11100011;
DRAM[56366] = 8'b11011111;
DRAM[56367] = 8'b11011101;
DRAM[56368] = 8'b11011101;
DRAM[56369] = 8'b11011011;
DRAM[56370] = 8'b11011001;
DRAM[56371] = 8'b11010111;
DRAM[56372] = 8'b11010110;
DRAM[56373] = 8'b11010011;
DRAM[56374] = 8'b11001110;
DRAM[56375] = 8'b11001011;
DRAM[56376] = 8'b11000111;
DRAM[56377] = 8'b11000101;
DRAM[56378] = 8'b11000010;
DRAM[56379] = 8'b11000000;
DRAM[56380] = 8'b10111111;
DRAM[56381] = 8'b10111110;
DRAM[56382] = 8'b10111011;
DRAM[56383] = 8'b10111001;
DRAM[56384] = 8'b10110010;
DRAM[56385] = 8'b10110000;
DRAM[56386] = 8'b10110110;
DRAM[56387] = 8'b10100110;
DRAM[56388] = 8'b10100010;
DRAM[56389] = 8'b10101011;
DRAM[56390] = 8'b10100011;
DRAM[56391] = 8'b10100011;
DRAM[56392] = 8'b10001001;
DRAM[56393] = 8'b10010111;
DRAM[56394] = 8'b10011001;
DRAM[56395] = 8'b10011101;
DRAM[56396] = 8'b10100111;
DRAM[56397] = 8'b10011011;
DRAM[56398] = 8'b10010000;
DRAM[56399] = 8'b10011101;
DRAM[56400] = 8'b10010101;
DRAM[56401] = 8'b10100100;
DRAM[56402] = 8'b10100000;
DRAM[56403] = 8'b10010010;
DRAM[56404] = 8'b10010011;
DRAM[56405] = 8'b10010100;
DRAM[56406] = 8'b10001100;
DRAM[56407] = 8'b10000111;
DRAM[56408] = 8'b10010001;
DRAM[56409] = 8'b10010000;
DRAM[56410] = 8'b10001111;
DRAM[56411] = 8'b10001000;
DRAM[56412] = 8'b10001001;
DRAM[56413] = 8'b10001001;
DRAM[56414] = 8'b10001000;
DRAM[56415] = 8'b10000010;
DRAM[56416] = 8'b1111011;
DRAM[56417] = 8'b1111100;
DRAM[56418] = 8'b1111010;
DRAM[56419] = 8'b1111010;
DRAM[56420] = 8'b1111101;
DRAM[56421] = 8'b1111110;
DRAM[56422] = 8'b1111111;
DRAM[56423] = 8'b10000101;
DRAM[56424] = 8'b1101111;
DRAM[56425] = 8'b1101101;
DRAM[56426] = 8'b1101011;
DRAM[56427] = 8'b1101010;
DRAM[56428] = 8'b1100110;
DRAM[56429] = 8'b1100000;
DRAM[56430] = 8'b1011110;
DRAM[56431] = 8'b1100000;
DRAM[56432] = 8'b1011010;
DRAM[56433] = 8'b1011110;
DRAM[56434] = 8'b1100011;
DRAM[56435] = 8'b1100101;
DRAM[56436] = 8'b1011110;
DRAM[56437] = 8'b1010101;
DRAM[56438] = 8'b1010000;
DRAM[56439] = 8'b1010001;
DRAM[56440] = 8'b1010011;
DRAM[56441] = 8'b1101010;
DRAM[56442] = 8'b1100000;
DRAM[56443] = 8'b1101100;
DRAM[56444] = 8'b1110001;
DRAM[56445] = 8'b1100011;
DRAM[56446] = 8'b1110010;
DRAM[56447] = 8'b1110011;
DRAM[56448] = 8'b1101101;
DRAM[56449] = 8'b1100011;
DRAM[56450] = 8'b1101000;
DRAM[56451] = 8'b1100001;
DRAM[56452] = 8'b1100000;
DRAM[56453] = 8'b1100100;
DRAM[56454] = 8'b1011001;
DRAM[56455] = 8'b1011110;
DRAM[56456] = 8'b1001101;
DRAM[56457] = 8'b1010100;
DRAM[56458] = 8'b1011101;
DRAM[56459] = 8'b1100000;
DRAM[56460] = 8'b1011000;
DRAM[56461] = 8'b1001110;
DRAM[56462] = 8'b1001110;
DRAM[56463] = 8'b1010101;
DRAM[56464] = 8'b1011101;
DRAM[56465] = 8'b1100011;
DRAM[56466] = 8'b1100001;
DRAM[56467] = 8'b1011010;
DRAM[56468] = 8'b1011011;
DRAM[56469] = 8'b1100101;
DRAM[56470] = 8'b1100101;
DRAM[56471] = 8'b1011100;
DRAM[56472] = 8'b1110000;
DRAM[56473] = 8'b1110001;
DRAM[56474] = 8'b1110100;
DRAM[56475] = 8'b1110111;
DRAM[56476] = 8'b1111100;
DRAM[56477] = 8'b10000000;
DRAM[56478] = 8'b10000000;
DRAM[56479] = 8'b1111110;
DRAM[56480] = 8'b1111110;
DRAM[56481] = 8'b1111111;
DRAM[56482] = 8'b10000010;
DRAM[56483] = 8'b10000110;
DRAM[56484] = 8'b10001100;
DRAM[56485] = 8'b10010011;
DRAM[56486] = 8'b10010111;
DRAM[56487] = 8'b10011001;
DRAM[56488] = 8'b10011110;
DRAM[56489] = 8'b10011100;
DRAM[56490] = 8'b10011110;
DRAM[56491] = 8'b10100101;
DRAM[56492] = 8'b10101101;
DRAM[56493] = 8'b10110000;
DRAM[56494] = 8'b10101100;
DRAM[56495] = 8'b10100110;
DRAM[56496] = 8'b10101101;
DRAM[56497] = 8'b10110000;
DRAM[56498] = 8'b10110100;
DRAM[56499] = 8'b10111001;
DRAM[56500] = 8'b10111101;
DRAM[56501] = 8'b10111111;
DRAM[56502] = 8'b10111110;
DRAM[56503] = 8'b10111101;
DRAM[56504] = 8'b11000011;
DRAM[56505] = 8'b11001000;
DRAM[56506] = 8'b11010001;
DRAM[56507] = 8'b11011111;
DRAM[56508] = 8'b11101100;
DRAM[56509] = 8'b11110101;
DRAM[56510] = 8'b11111001;
DRAM[56511] = 8'b11111001;
DRAM[56512] = 8'b11101110;
DRAM[56513] = 8'b11110000;
DRAM[56514] = 8'b11101001;
DRAM[56515] = 8'b11010010;
DRAM[56516] = 8'b10110100;
DRAM[56517] = 8'b10011100;
DRAM[56518] = 8'b10010000;
DRAM[56519] = 8'b10001100;
DRAM[56520] = 8'b10000111;
DRAM[56521] = 8'b10000111;
DRAM[56522] = 8'b10000111;
DRAM[56523] = 8'b10000110;
DRAM[56524] = 8'b10000110;
DRAM[56525] = 8'b10000101;
DRAM[56526] = 8'b10000101;
DRAM[56527] = 8'b10000100;
DRAM[56528] = 8'b1111111;
DRAM[56529] = 8'b1111110;
DRAM[56530] = 8'b1111100;
DRAM[56531] = 8'b1111011;
DRAM[56532] = 8'b1111001;
DRAM[56533] = 8'b1111000;
DRAM[56534] = 8'b1111000;
DRAM[56535] = 8'b1111000;
DRAM[56536] = 8'b1111000;
DRAM[56537] = 8'b1110110;
DRAM[56538] = 8'b1110011;
DRAM[56539] = 8'b1110010;
DRAM[56540] = 8'b1110010;
DRAM[56541] = 8'b1110001;
DRAM[56542] = 8'b1101111;
DRAM[56543] = 8'b1101101;
DRAM[56544] = 8'b1101111;
DRAM[56545] = 8'b1101110;
DRAM[56546] = 8'b1101101;
DRAM[56547] = 8'b1101100;
DRAM[56548] = 8'b1101100;
DRAM[56549] = 8'b1101100;
DRAM[56550] = 8'b1101100;
DRAM[56551] = 8'b1101100;
DRAM[56552] = 8'b1101011;
DRAM[56553] = 8'b1101011;
DRAM[56554] = 8'b1101010;
DRAM[56555] = 8'b1101001;
DRAM[56556] = 8'b1101000;
DRAM[56557] = 8'b1101001;
DRAM[56558] = 8'b1101001;
DRAM[56559] = 8'b1101001;
DRAM[56560] = 8'b1101011;
DRAM[56561] = 8'b1101011;
DRAM[56562] = 8'b1101010;
DRAM[56563] = 8'b1101010;
DRAM[56564] = 8'b1101010;
DRAM[56565] = 8'b1101010;
DRAM[56566] = 8'b1101001;
DRAM[56567] = 8'b1101001;
DRAM[56568] = 8'b1101001;
DRAM[56569] = 8'b1101001;
DRAM[56570] = 8'b1101010;
DRAM[56571] = 8'b1101010;
DRAM[56572] = 8'b1101010;
DRAM[56573] = 8'b1101010;
DRAM[56574] = 8'b1101011;
DRAM[56575] = 8'b1101011;
DRAM[56576] = 8'b10001101;
DRAM[56577] = 8'b10001110;
DRAM[56578] = 8'b10001111;
DRAM[56579] = 8'b10010001;
DRAM[56580] = 8'b10010010;
DRAM[56581] = 8'b10010100;
DRAM[56582] = 8'b10010101;
DRAM[56583] = 8'b10010110;
DRAM[56584] = 8'b10011000;
DRAM[56585] = 8'b10011010;
DRAM[56586] = 8'b10011101;
DRAM[56587] = 8'b10011110;
DRAM[56588] = 8'b10011110;
DRAM[56589] = 8'b10011111;
DRAM[56590] = 8'b10100010;
DRAM[56591] = 8'b10100100;
DRAM[56592] = 8'b10101110;
DRAM[56593] = 8'b10111110;
DRAM[56594] = 8'b11010110;
DRAM[56595] = 8'b11101011;
DRAM[56596] = 8'b11111000;
DRAM[56597] = 8'b11111100;
DRAM[56598] = 8'b11111100;
DRAM[56599] = 8'b11111010;
DRAM[56600] = 8'b11111101;
DRAM[56601] = 8'b11111100;
DRAM[56602] = 8'b11111011;
DRAM[56603] = 8'b11111010;
DRAM[56604] = 8'b11110111;
DRAM[56605] = 8'b11110101;
DRAM[56606] = 8'b11110010;
DRAM[56607] = 8'b11110001;
DRAM[56608] = 8'b11100101;
DRAM[56609] = 8'b11101001;
DRAM[56610] = 8'b11101110;
DRAM[56611] = 8'b11110010;
DRAM[56612] = 8'b11110011;
DRAM[56613] = 8'b11110001;
DRAM[56614] = 8'b11101110;
DRAM[56615] = 8'b11101100;
DRAM[56616] = 8'b11110111;
DRAM[56617] = 8'b11110001;
DRAM[56618] = 8'b11101000;
DRAM[56619] = 8'b11100011;
DRAM[56620] = 8'b11100001;
DRAM[56621] = 8'b11100010;
DRAM[56622] = 8'b11100011;
DRAM[56623] = 8'b11100011;
DRAM[56624] = 8'b11011111;
DRAM[56625] = 8'b11011011;
DRAM[56626] = 8'b11010111;
DRAM[56627] = 8'b11010100;
DRAM[56628] = 8'b11010011;
DRAM[56629] = 8'b11010010;
DRAM[56630] = 8'b11010000;
DRAM[56631] = 8'b11001111;
DRAM[56632] = 8'b11001110;
DRAM[56633] = 8'b11001011;
DRAM[56634] = 8'b11001000;
DRAM[56635] = 8'b11000110;
DRAM[56636] = 8'b11000100;
DRAM[56637] = 8'b11000000;
DRAM[56638] = 8'b10111100;
DRAM[56639] = 8'b10111000;
DRAM[56640] = 8'b10100001;
DRAM[56641] = 8'b10101011;
DRAM[56642] = 8'b10111001;
DRAM[56643] = 8'b10101011;
DRAM[56644] = 8'b10101000;
DRAM[56645] = 8'b10110000;
DRAM[56646] = 8'b10011001;
DRAM[56647] = 8'b10001001;
DRAM[56648] = 8'b10001011;
DRAM[56649] = 8'b10001100;
DRAM[56650] = 8'b10001100;
DRAM[56651] = 8'b10010011;
DRAM[56652] = 8'b10011010;
DRAM[56653] = 8'b10010110;
DRAM[56654] = 8'b10010111;
DRAM[56655] = 8'b10100101;
DRAM[56656] = 8'b10010110;
DRAM[56657] = 8'b10010100;
DRAM[56658] = 8'b10010000;
DRAM[56659] = 8'b10010110;
DRAM[56660] = 8'b10011001;
DRAM[56661] = 8'b10001100;
DRAM[56662] = 8'b10000110;
DRAM[56663] = 8'b10010011;
DRAM[56664] = 8'b10010011;
DRAM[56665] = 8'b10010000;
DRAM[56666] = 8'b10010010;
DRAM[56667] = 8'b10000111;
DRAM[56668] = 8'b10001110;
DRAM[56669] = 8'b10001001;
DRAM[56670] = 8'b10001101;
DRAM[56671] = 8'b10000101;
DRAM[56672] = 8'b1111100;
DRAM[56673] = 8'b10000011;
DRAM[56674] = 8'b1111101;
DRAM[56675] = 8'b1111000;
DRAM[56676] = 8'b1111111;
DRAM[56677] = 8'b10000000;
DRAM[56678] = 8'b1111101;
DRAM[56679] = 8'b10000001;
DRAM[56680] = 8'b1110000;
DRAM[56681] = 8'b1101110;
DRAM[56682] = 8'b1101100;
DRAM[56683] = 8'b1101001;
DRAM[56684] = 8'b1100110;
DRAM[56685] = 8'b1100010;
DRAM[56686] = 8'b1100000;
DRAM[56687] = 8'b1011111;
DRAM[56688] = 8'b1011101;
DRAM[56689] = 8'b1100001;
DRAM[56690] = 8'b1100110;
DRAM[56691] = 8'b1100101;
DRAM[56692] = 8'b1011111;
DRAM[56693] = 8'b1010111;
DRAM[56694] = 8'b1010010;
DRAM[56695] = 8'b1010001;
DRAM[56696] = 8'b1010010;
DRAM[56697] = 8'b1100100;
DRAM[56698] = 8'b1100101;
DRAM[56699] = 8'b1101101;
DRAM[56700] = 8'b1110000;
DRAM[56701] = 8'b1100110;
DRAM[56702] = 8'b1101101;
DRAM[56703] = 8'b1111000;
DRAM[56704] = 8'b1110001;
DRAM[56705] = 8'b1100100;
DRAM[56706] = 8'b1100111;
DRAM[56707] = 8'b1100000;
DRAM[56708] = 8'b1011111;
DRAM[56709] = 8'b1100011;
DRAM[56710] = 8'b1011011;
DRAM[56711] = 8'b1100100;
DRAM[56712] = 8'b1001111;
DRAM[56713] = 8'b1010100;
DRAM[56714] = 8'b1011101;
DRAM[56715] = 8'b1100011;
DRAM[56716] = 8'b1100000;
DRAM[56717] = 8'b1011000;
DRAM[56718] = 8'b1010110;
DRAM[56719] = 8'b1011010;
DRAM[56720] = 8'b1011000;
DRAM[56721] = 8'b1100101;
DRAM[56722] = 8'b1100101;
DRAM[56723] = 8'b1011010;
DRAM[56724] = 8'b1011011;
DRAM[56725] = 8'b1101000;
DRAM[56726] = 8'b1101010;
DRAM[56727] = 8'b1011111;
DRAM[56728] = 8'b1101110;
DRAM[56729] = 8'b1110010;
DRAM[56730] = 8'b1110101;
DRAM[56731] = 8'b1110101;
DRAM[56732] = 8'b1111001;
DRAM[56733] = 8'b1111110;
DRAM[56734] = 8'b10000001;
DRAM[56735] = 8'b10000000;
DRAM[56736] = 8'b10000010;
DRAM[56737] = 8'b10000000;
DRAM[56738] = 8'b1111110;
DRAM[56739] = 8'b10000001;
DRAM[56740] = 8'b10000111;
DRAM[56741] = 8'b10001110;
DRAM[56742] = 8'b10010100;
DRAM[56743] = 8'b10010111;
DRAM[56744] = 8'b10011001;
DRAM[56745] = 8'b10011111;
DRAM[56746] = 8'b10100100;
DRAM[56747] = 8'b10100101;
DRAM[56748] = 8'b10100100;
DRAM[56749] = 8'b10101000;
DRAM[56750] = 8'b10110001;
DRAM[56751] = 8'b10111001;
DRAM[56752] = 8'b10110010;
DRAM[56753] = 8'b10110010;
DRAM[56754] = 8'b10110101;
DRAM[56755] = 8'b10111001;
DRAM[56756] = 8'b10111110;
DRAM[56757] = 8'b11000000;
DRAM[56758] = 8'b11000000;
DRAM[56759] = 8'b10111111;
DRAM[56760] = 8'b11001010;
DRAM[56761] = 8'b11001100;
DRAM[56762] = 8'b11010010;
DRAM[56763] = 8'b11011110;
DRAM[56764] = 8'b11101100;
DRAM[56765] = 8'b11110110;
DRAM[56766] = 8'b11111000;
DRAM[56767] = 8'b11110111;
DRAM[56768] = 8'b11111101;
DRAM[56769] = 8'b11100100;
DRAM[56770] = 8'b11000011;
DRAM[56771] = 8'b10110001;
DRAM[56772] = 8'b10101111;
DRAM[56773] = 8'b10101101;
DRAM[56774] = 8'b10011100;
DRAM[56775] = 8'b10001001;
DRAM[56776] = 8'b10001011;
DRAM[56777] = 8'b10001001;
DRAM[56778] = 8'b10000111;
DRAM[56779] = 8'b10000101;
DRAM[56780] = 8'b10000100;
DRAM[56781] = 8'b10000100;
DRAM[56782] = 8'b10000101;
DRAM[56783] = 8'b10000110;
DRAM[56784] = 8'b10000001;
DRAM[56785] = 8'b10000000;
DRAM[56786] = 8'b1111110;
DRAM[56787] = 8'b1111011;
DRAM[56788] = 8'b1111001;
DRAM[56789] = 8'b1111000;
DRAM[56790] = 8'b1110111;
DRAM[56791] = 8'b1110111;
DRAM[56792] = 8'b1110111;
DRAM[56793] = 8'b1110101;
DRAM[56794] = 8'b1110011;
DRAM[56795] = 8'b1110010;
DRAM[56796] = 8'b1110010;
DRAM[56797] = 8'b1110001;
DRAM[56798] = 8'b1101111;
DRAM[56799] = 8'b1101100;
DRAM[56800] = 8'b1101110;
DRAM[56801] = 8'b1101101;
DRAM[56802] = 8'b1101100;
DRAM[56803] = 8'b1101100;
DRAM[56804] = 8'b1101011;
DRAM[56805] = 8'b1101100;
DRAM[56806] = 8'b1101100;
DRAM[56807] = 8'b1101101;
DRAM[56808] = 8'b1101011;
DRAM[56809] = 8'b1101011;
DRAM[56810] = 8'b1101010;
DRAM[56811] = 8'b1101001;
DRAM[56812] = 8'b1101000;
DRAM[56813] = 8'b1101000;
DRAM[56814] = 8'b1101001;
DRAM[56815] = 8'b1101001;
DRAM[56816] = 8'b1101010;
DRAM[56817] = 8'b1101010;
DRAM[56818] = 8'b1101010;
DRAM[56819] = 8'b1101010;
DRAM[56820] = 8'b1101010;
DRAM[56821] = 8'b1101010;
DRAM[56822] = 8'b1101010;
DRAM[56823] = 8'b1101010;
DRAM[56824] = 8'b1101010;
DRAM[56825] = 8'b1101010;
DRAM[56826] = 8'b1101010;
DRAM[56827] = 8'b1101010;
DRAM[56828] = 8'b1101010;
DRAM[56829] = 8'b1101010;
DRAM[56830] = 8'b1101010;
DRAM[56831] = 8'b1101010;
DRAM[56832] = 8'b10001100;
DRAM[56833] = 8'b10001101;
DRAM[56834] = 8'b10001110;
DRAM[56835] = 8'b10010000;
DRAM[56836] = 8'b10010001;
DRAM[56837] = 8'b10010011;
DRAM[56838] = 8'b10010100;
DRAM[56839] = 8'b10010101;
DRAM[56840] = 8'b10010110;
DRAM[56841] = 8'b10011000;
DRAM[56842] = 8'b10011011;
DRAM[56843] = 8'b10011100;
DRAM[56844] = 8'b10011101;
DRAM[56845] = 8'b10011110;
DRAM[56846] = 8'b10100001;
DRAM[56847] = 8'b10100011;
DRAM[56848] = 8'b10110000;
DRAM[56849] = 8'b11000011;
DRAM[56850] = 8'b11011110;
DRAM[56851] = 8'b11110001;
DRAM[56852] = 8'b11111001;
DRAM[56853] = 8'b11111010;
DRAM[56854] = 8'b11111100;
DRAM[56855] = 8'b11111101;
DRAM[56856] = 8'b11111100;
DRAM[56857] = 8'b11111011;
DRAM[56858] = 8'b11111010;
DRAM[56859] = 8'b11111000;
DRAM[56860] = 8'b11110101;
DRAM[56861] = 8'b11110010;
DRAM[56862] = 8'b11110000;
DRAM[56863] = 8'b11101110;
DRAM[56864] = 8'b11100011;
DRAM[56865] = 8'b11101001;
DRAM[56866] = 8'b11101110;
DRAM[56867] = 8'b11101111;
DRAM[56868] = 8'b11101110;
DRAM[56869] = 8'b11101101;
DRAM[56870] = 8'b11101111;
DRAM[56871] = 8'b11110010;
DRAM[56872] = 8'b11101100;
DRAM[56873] = 8'b11100110;
DRAM[56874] = 8'b11100000;
DRAM[56875] = 8'b11011111;
DRAM[56876] = 8'b11100011;
DRAM[56877] = 8'b11100111;
DRAM[56878] = 8'b11100110;
DRAM[56879] = 8'b11100100;
DRAM[56880] = 8'b11011001;
DRAM[56881] = 8'b11010111;
DRAM[56882] = 8'b11010101;
DRAM[56883] = 8'b11010011;
DRAM[56884] = 8'b11010011;
DRAM[56885] = 8'b11010001;
DRAM[56886] = 8'b11001110;
DRAM[56887] = 8'b11001100;
DRAM[56888] = 8'b11000110;
DRAM[56889] = 8'b11000011;
DRAM[56890] = 8'b10111110;
DRAM[56891] = 8'b10111011;
DRAM[56892] = 8'b10111001;
DRAM[56893] = 8'b10111000;
DRAM[56894] = 8'b10110101;
DRAM[56895] = 8'b10110011;
DRAM[56896] = 8'b10110010;
DRAM[56897] = 8'b10101010;
DRAM[56898] = 8'b10101001;
DRAM[56899] = 8'b10011010;
DRAM[56900] = 8'b10011011;
DRAM[56901] = 8'b10100111;
DRAM[56902] = 8'b10011011;
DRAM[56903] = 8'b10010111;
DRAM[56904] = 8'b10010101;
DRAM[56905] = 8'b10001000;
DRAM[56906] = 8'b10001010;
DRAM[56907] = 8'b10010100;
DRAM[56908] = 8'b10010100;
DRAM[56909] = 8'b10010101;
DRAM[56910] = 8'b10011101;
DRAM[56911] = 8'b10100001;
DRAM[56912] = 8'b10001100;
DRAM[56913] = 8'b10001110;
DRAM[56914] = 8'b10001111;
DRAM[56915] = 8'b10010101;
DRAM[56916] = 8'b10010111;
DRAM[56917] = 8'b10001010;
DRAM[56918] = 8'b10001001;
DRAM[56919] = 8'b10011011;
DRAM[56920] = 8'b10010111;
DRAM[56921] = 8'b10010100;
DRAM[56922] = 8'b10011010;
DRAM[56923] = 8'b10001100;
DRAM[56924] = 8'b10010110;
DRAM[56925] = 8'b10001011;
DRAM[56926] = 8'b10001111;
DRAM[56927] = 8'b10000100;
DRAM[56928] = 8'b1111110;
DRAM[56929] = 8'b10001001;
DRAM[56930] = 8'b1111111;
DRAM[56931] = 8'b1110101;
DRAM[56932] = 8'b10000000;
DRAM[56933] = 8'b10000010;
DRAM[56934] = 8'b1111001;
DRAM[56935] = 8'b1111100;
DRAM[56936] = 8'b1110011;
DRAM[56937] = 8'b1110010;
DRAM[56938] = 8'b1101111;
DRAM[56939] = 8'b1101011;
DRAM[56940] = 8'b1101001;
DRAM[56941] = 8'b1100111;
DRAM[56942] = 8'b1100100;
DRAM[56943] = 8'b1100001;
DRAM[56944] = 8'b1100000;
DRAM[56945] = 8'b1100011;
DRAM[56946] = 8'b1100110;
DRAM[56947] = 8'b1100101;
DRAM[56948] = 8'b1100010;
DRAM[56949] = 8'b1011101;
DRAM[56950] = 8'b1011000;
DRAM[56951] = 8'b1010100;
DRAM[56952] = 8'b1010110;
DRAM[56953] = 8'b1011010;
DRAM[56954] = 8'b1100110;
DRAM[56955] = 8'b1101000;
DRAM[56956] = 8'b1101110;
DRAM[56957] = 8'b1101101;
DRAM[56958] = 8'b1100110;
DRAM[56959] = 8'b1110111;
DRAM[56960] = 8'b1110101;
DRAM[56961] = 8'b1100101;
DRAM[56962] = 8'b1100111;
DRAM[56963] = 8'b1100000;
DRAM[56964] = 8'b1100000;
DRAM[56965] = 8'b1100110;
DRAM[56966] = 8'b1100001;
DRAM[56967] = 8'b1101100;
DRAM[56968] = 8'b1011011;
DRAM[56969] = 8'b1011010;
DRAM[56970] = 8'b1011110;
DRAM[56971] = 8'b1100101;
DRAM[56972] = 8'b1101000;
DRAM[56973] = 8'b1100100;
DRAM[56974] = 8'b1100001;
DRAM[56975] = 8'b1100001;
DRAM[56976] = 8'b1011011;
DRAM[56977] = 8'b1100100;
DRAM[56978] = 8'b1101001;
DRAM[56979] = 8'b1100101;
DRAM[56980] = 8'b1100011;
DRAM[56981] = 8'b1100111;
DRAM[56982] = 8'b1101000;
DRAM[56983] = 8'b1100101;
DRAM[56984] = 8'b1100101;
DRAM[56985] = 8'b1101110;
DRAM[56986] = 8'b1110101;
DRAM[56987] = 8'b1110110;
DRAM[56988] = 8'b1111001;
DRAM[56989] = 8'b10000000;
DRAM[56990] = 8'b10000101;
DRAM[56991] = 8'b10000101;
DRAM[56992] = 8'b10001001;
DRAM[56993] = 8'b10000101;
DRAM[56994] = 8'b10000010;
DRAM[56995] = 8'b10000011;
DRAM[56996] = 8'b10001000;
DRAM[56997] = 8'b10001110;
DRAM[56998] = 8'b10010011;
DRAM[56999] = 8'b10010100;
DRAM[57000] = 8'b10010110;
DRAM[57001] = 8'b10011011;
DRAM[57002] = 8'b10100001;
DRAM[57003] = 8'b10100010;
DRAM[57004] = 8'b10100010;
DRAM[57005] = 8'b10100101;
DRAM[57006] = 8'b10101101;
DRAM[57007] = 8'b10110101;
DRAM[57008] = 8'b10110010;
DRAM[57009] = 8'b10110001;
DRAM[57010] = 8'b10110001;
DRAM[57011] = 8'b10110101;
DRAM[57012] = 8'b10111011;
DRAM[57013] = 8'b11000000;
DRAM[57014] = 8'b11000010;
DRAM[57015] = 8'b11000010;
DRAM[57016] = 8'b11001000;
DRAM[57017] = 8'b11001101;
DRAM[57018] = 8'b11010110;
DRAM[57019] = 8'b11100001;
DRAM[57020] = 8'b11101100;
DRAM[57021] = 8'b11110011;
DRAM[57022] = 8'b11110111;
DRAM[57023] = 8'b11111000;
DRAM[57024] = 8'b11111111;
DRAM[57025] = 8'b11110110;
DRAM[57026] = 8'b11010110;
DRAM[57027] = 8'b10101010;
DRAM[57028] = 8'b10001010;
DRAM[57029] = 8'b10000001;
DRAM[57030] = 8'b10001000;
DRAM[57031] = 8'b10001110;
DRAM[57032] = 8'b10001010;
DRAM[57033] = 8'b10001001;
DRAM[57034] = 8'b10000111;
DRAM[57035] = 8'b10000110;
DRAM[57036] = 8'b10000101;
DRAM[57037] = 8'b10000101;
DRAM[57038] = 8'b10000101;
DRAM[57039] = 8'b10000101;
DRAM[57040] = 8'b1111111;
DRAM[57041] = 8'b1111110;
DRAM[57042] = 8'b1111100;
DRAM[57043] = 8'b1111010;
DRAM[57044] = 8'b1111001;
DRAM[57045] = 8'b1111000;
DRAM[57046] = 8'b1110111;
DRAM[57047] = 8'b1110111;
DRAM[57048] = 8'b1111000;
DRAM[57049] = 8'b1110110;
DRAM[57050] = 8'b1110100;
DRAM[57051] = 8'b1110011;
DRAM[57052] = 8'b1110011;
DRAM[57053] = 8'b1110010;
DRAM[57054] = 8'b1101111;
DRAM[57055] = 8'b1101101;
DRAM[57056] = 8'b1101100;
DRAM[57057] = 8'b1101100;
DRAM[57058] = 8'b1101011;
DRAM[57059] = 8'b1101011;
DRAM[57060] = 8'b1101011;
DRAM[57061] = 8'b1101100;
DRAM[57062] = 8'b1101101;
DRAM[57063] = 8'b1101110;
DRAM[57064] = 8'b1101100;
DRAM[57065] = 8'b1101011;
DRAM[57066] = 8'b1101010;
DRAM[57067] = 8'b1101001;
DRAM[57068] = 8'b1101001;
DRAM[57069] = 8'b1101001;
DRAM[57070] = 8'b1101001;
DRAM[57071] = 8'b1101001;
DRAM[57072] = 8'b1101010;
DRAM[57073] = 8'b1101010;
DRAM[57074] = 8'b1101010;
DRAM[57075] = 8'b1101010;
DRAM[57076] = 8'b1101010;
DRAM[57077] = 8'b1101010;
DRAM[57078] = 8'b1101010;
DRAM[57079] = 8'b1101010;
DRAM[57080] = 8'b1101010;
DRAM[57081] = 8'b1101010;
DRAM[57082] = 8'b1101010;
DRAM[57083] = 8'b1101010;
DRAM[57084] = 8'b1101010;
DRAM[57085] = 8'b1101010;
DRAM[57086] = 8'b1101010;
DRAM[57087] = 8'b1101010;
DRAM[57088] = 8'b10001100;
DRAM[57089] = 8'b10001100;
DRAM[57090] = 8'b10001101;
DRAM[57091] = 8'b10001111;
DRAM[57092] = 8'b10010001;
DRAM[57093] = 8'b10010010;
DRAM[57094] = 8'b10010011;
DRAM[57095] = 8'b10010100;
DRAM[57096] = 8'b10010101;
DRAM[57097] = 8'b10010111;
DRAM[57098] = 8'b10011010;
DRAM[57099] = 8'b10011011;
DRAM[57100] = 8'b10011100;
DRAM[57101] = 8'b10011110;
DRAM[57102] = 8'b10100001;
DRAM[57103] = 8'b10100011;
DRAM[57104] = 8'b10110001;
DRAM[57105] = 8'b11000111;
DRAM[57106] = 8'b11100011;
DRAM[57107] = 8'b11110100;
DRAM[57108] = 8'b11111001;
DRAM[57109] = 8'b11111001;
DRAM[57110] = 8'b11111100;
DRAM[57111] = 8'b11111111;
DRAM[57112] = 8'b11111011;
DRAM[57113] = 8'b11111010;
DRAM[57114] = 8'b11111001;
DRAM[57115] = 8'b11110111;
DRAM[57116] = 8'b11110100;
DRAM[57117] = 8'b11110001;
DRAM[57118] = 8'b11101110;
DRAM[57119] = 8'b11101101;
DRAM[57120] = 8'b11101100;
DRAM[57121] = 8'b11110000;
DRAM[57122] = 8'b11110010;
DRAM[57123] = 8'b11101111;
DRAM[57124] = 8'b11101000;
DRAM[57125] = 8'b11100110;
DRAM[57126] = 8'b11101011;
DRAM[57127] = 8'b11110001;
DRAM[57128] = 8'b11100111;
DRAM[57129] = 8'b11100100;
DRAM[57130] = 8'b11100100;
DRAM[57131] = 8'b11101001;
DRAM[57132] = 8'b11101110;
DRAM[57133] = 8'b11101101;
DRAM[57134] = 8'b11100100;
DRAM[57135] = 8'b11011011;
DRAM[57136] = 8'b11011100;
DRAM[57137] = 8'b11011011;
DRAM[57138] = 8'b11011001;
DRAM[57139] = 8'b11010110;
DRAM[57140] = 8'b11010001;
DRAM[57141] = 8'b11001010;
DRAM[57142] = 8'b11000001;
DRAM[57143] = 8'b10111011;
DRAM[57144] = 8'b10110111;
DRAM[57145] = 8'b10110011;
DRAM[57146] = 8'b10101101;
DRAM[57147] = 8'b10101001;
DRAM[57148] = 8'b10101001;
DRAM[57149] = 8'b10101010;
DRAM[57150] = 8'b10101010;
DRAM[57151] = 8'b10101010;
DRAM[57152] = 8'b10100001;
DRAM[57153] = 8'b10010110;
DRAM[57154] = 8'b10011111;
DRAM[57155] = 8'b10100010;
DRAM[57156] = 8'b10100111;
DRAM[57157] = 8'b10100110;
DRAM[57158] = 8'b10001111;
DRAM[57159] = 8'b10001011;
DRAM[57160] = 8'b10011110;
DRAM[57161] = 8'b10001010;
DRAM[57162] = 8'b10010001;
DRAM[57163] = 8'b10011111;
DRAM[57164] = 8'b10011000;
DRAM[57165] = 8'b10010110;
DRAM[57166] = 8'b10011100;
DRAM[57167] = 8'b10010111;
DRAM[57168] = 8'b10001100;
DRAM[57169] = 8'b10100011;
DRAM[57170] = 8'b10100100;
DRAM[57171] = 8'b10010101;
DRAM[57172] = 8'b10001111;
DRAM[57173] = 8'b10001111;
DRAM[57174] = 8'b10010000;
DRAM[57175] = 8'b10010100;
DRAM[57176] = 8'b10010100;
DRAM[57177] = 8'b10010010;
DRAM[57178] = 8'b10011011;
DRAM[57179] = 8'b10001011;
DRAM[57180] = 8'b10010111;
DRAM[57181] = 8'b10000111;
DRAM[57182] = 8'b10001001;
DRAM[57183] = 8'b1111100;
DRAM[57184] = 8'b10000001;
DRAM[57185] = 8'b10001101;
DRAM[57186] = 8'b10000000;
DRAM[57187] = 8'b1110101;
DRAM[57188] = 8'b10000010;
DRAM[57189] = 8'b10000100;
DRAM[57190] = 8'b1111000;
DRAM[57191] = 8'b1111010;
DRAM[57192] = 8'b1111000;
DRAM[57193] = 8'b1110111;
DRAM[57194] = 8'b1110011;
DRAM[57195] = 8'b1101111;
DRAM[57196] = 8'b1101101;
DRAM[57197] = 8'b1101011;
DRAM[57198] = 8'b1101000;
DRAM[57199] = 8'b1100100;
DRAM[57200] = 8'b1100001;
DRAM[57201] = 8'b1100100;
DRAM[57202] = 8'b1100110;
DRAM[57203] = 8'b1100101;
DRAM[57204] = 8'b1100100;
DRAM[57205] = 8'b1100001;
DRAM[57206] = 8'b1011101;
DRAM[57207] = 8'b1011000;
DRAM[57208] = 8'b1011001;
DRAM[57209] = 8'b1010011;
DRAM[57210] = 8'b1100100;
DRAM[57211] = 8'b1100011;
DRAM[57212] = 8'b1101101;
DRAM[57213] = 8'b1110011;
DRAM[57214] = 8'b1100000;
DRAM[57215] = 8'b1110011;
DRAM[57216] = 8'b1111001;
DRAM[57217] = 8'b1101000;
DRAM[57218] = 8'b1101001;
DRAM[57219] = 8'b1100010;
DRAM[57220] = 8'b1100011;
DRAM[57221] = 8'b1101010;
DRAM[57222] = 8'b1100111;
DRAM[57223] = 8'b1110100;
DRAM[57224] = 8'b1100101;
DRAM[57225] = 8'b1011110;
DRAM[57226] = 8'b1011100;
DRAM[57227] = 8'b1100010;
DRAM[57228] = 8'b1100110;
DRAM[57229] = 8'b1100101;
DRAM[57230] = 8'b1100001;
DRAM[57231] = 8'b1011111;
DRAM[57232] = 8'b1100011;
DRAM[57233] = 8'b1100101;
DRAM[57234] = 8'b1101100;
DRAM[57235] = 8'b1110010;
DRAM[57236] = 8'b1101100;
DRAM[57237] = 8'b1100010;
DRAM[57238] = 8'b1100001;
DRAM[57239] = 8'b1100110;
DRAM[57240] = 8'b1011001;
DRAM[57241] = 8'b1100111;
DRAM[57242] = 8'b1110100;
DRAM[57243] = 8'b1111000;
DRAM[57244] = 8'b1111011;
DRAM[57245] = 8'b10000100;
DRAM[57246] = 8'b10001010;
DRAM[57247] = 8'b10001011;
DRAM[57248] = 8'b10001111;
DRAM[57249] = 8'b10001011;
DRAM[57250] = 8'b10001000;
DRAM[57251] = 8'b10001000;
DRAM[57252] = 8'b10001101;
DRAM[57253] = 8'b10010010;
DRAM[57254] = 8'b10010100;
DRAM[57255] = 8'b10010100;
DRAM[57256] = 8'b10010101;
DRAM[57257] = 8'b10010100;
DRAM[57258] = 8'b10010110;
DRAM[57259] = 8'b10011111;
DRAM[57260] = 8'b10101000;
DRAM[57261] = 8'b10101011;
DRAM[57262] = 8'b10100101;
DRAM[57263] = 8'b10011111;
DRAM[57264] = 8'b10101110;
DRAM[57265] = 8'b10101100;
DRAM[57266] = 8'b10101100;
DRAM[57267] = 8'b10110000;
DRAM[57268] = 8'b10111001;
DRAM[57269] = 8'b11000000;
DRAM[57270] = 8'b11000100;
DRAM[57271] = 8'b11000110;
DRAM[57272] = 8'b10111110;
DRAM[57273] = 8'b11001001;
DRAM[57274] = 8'b11010111;
DRAM[57275] = 8'b11100011;
DRAM[57276] = 8'b11101011;
DRAM[57277] = 8'b11110001;
DRAM[57278] = 8'b11110111;
DRAM[57279] = 8'b11111011;
DRAM[57280] = 8'b11110101;
DRAM[57281] = 8'b11101100;
DRAM[57282] = 8'b11010100;
DRAM[57283] = 8'b10110001;
DRAM[57284] = 8'b10011000;
DRAM[57285] = 8'b10001101;
DRAM[57286] = 8'b10001010;
DRAM[57287] = 8'b10000111;
DRAM[57288] = 8'b10000111;
DRAM[57289] = 8'b10000111;
DRAM[57290] = 8'b10000111;
DRAM[57291] = 8'b10000111;
DRAM[57292] = 8'b10000110;
DRAM[57293] = 8'b10000110;
DRAM[57294] = 8'b10000101;
DRAM[57295] = 8'b10000101;
DRAM[57296] = 8'b1111011;
DRAM[57297] = 8'b1111011;
DRAM[57298] = 8'b1111010;
DRAM[57299] = 8'b1111000;
DRAM[57300] = 8'b1111000;
DRAM[57301] = 8'b1111000;
DRAM[57302] = 8'b1111000;
DRAM[57303] = 8'b1111000;
DRAM[57304] = 8'b1111001;
DRAM[57305] = 8'b1110111;
DRAM[57306] = 8'b1110101;
DRAM[57307] = 8'b1110100;
DRAM[57308] = 8'b1110100;
DRAM[57309] = 8'b1110011;
DRAM[57310] = 8'b1110001;
DRAM[57311] = 8'b1101111;
DRAM[57312] = 8'b1101011;
DRAM[57313] = 8'b1101011;
DRAM[57314] = 8'b1101011;
DRAM[57315] = 8'b1101011;
DRAM[57316] = 8'b1101011;
DRAM[57317] = 8'b1101101;
DRAM[57318] = 8'b1101110;
DRAM[57319] = 8'b1101110;
DRAM[57320] = 8'b1101100;
DRAM[57321] = 8'b1101011;
DRAM[57322] = 8'b1101010;
DRAM[57323] = 8'b1101001;
DRAM[57324] = 8'b1101001;
DRAM[57325] = 8'b1101001;
DRAM[57326] = 8'b1101010;
DRAM[57327] = 8'b1101010;
DRAM[57328] = 8'b1101010;
DRAM[57329] = 8'b1101010;
DRAM[57330] = 8'b1101010;
DRAM[57331] = 8'b1101010;
DRAM[57332] = 8'b1101010;
DRAM[57333] = 8'b1101010;
DRAM[57334] = 8'b1101010;
DRAM[57335] = 8'b1101010;
DRAM[57336] = 8'b1101010;
DRAM[57337] = 8'b1101010;
DRAM[57338] = 8'b1101010;
DRAM[57339] = 8'b1101010;
DRAM[57340] = 8'b1101010;
DRAM[57341] = 8'b1101010;
DRAM[57342] = 8'b1101010;
DRAM[57343] = 8'b1101010;
DRAM[57344] = 8'b10010001;
DRAM[57345] = 8'b10001111;
DRAM[57346] = 8'b10001101;
DRAM[57347] = 8'b10001011;
DRAM[57348] = 8'b10001011;
DRAM[57349] = 8'b10001101;
DRAM[57350] = 8'b10010000;
DRAM[57351] = 8'b10010010;
DRAM[57352] = 8'b10011001;
DRAM[57353] = 8'b10010111;
DRAM[57354] = 8'b10011000;
DRAM[57355] = 8'b10011011;
DRAM[57356] = 8'b10011101;
DRAM[57357] = 8'b10011101;
DRAM[57358] = 8'b10100011;
DRAM[57359] = 8'b10101010;
DRAM[57360] = 8'b10111001;
DRAM[57361] = 8'b11010101;
DRAM[57362] = 8'b11101110;
DRAM[57363] = 8'b11110101;
DRAM[57364] = 8'b11110111;
DRAM[57365] = 8'b11111110;
DRAM[57366] = 8'b11111111;
DRAM[57367] = 8'b11111101;
DRAM[57368] = 8'b11111101;
DRAM[57369] = 8'b11111010;
DRAM[57370] = 8'b11110101;
DRAM[57371] = 8'b11110011;
DRAM[57372] = 8'b11110011;
DRAM[57373] = 8'b11110011;
DRAM[57374] = 8'b11110010;
DRAM[57375] = 8'b11110001;
DRAM[57376] = 8'b11101001;
DRAM[57377] = 8'b11101101;
DRAM[57378] = 8'b11110001;
DRAM[57379] = 8'b11110001;
DRAM[57380] = 8'b11101110;
DRAM[57381] = 8'b11101100;
DRAM[57382] = 8'b11101101;
DRAM[57383] = 8'b11101111;
DRAM[57384] = 8'b11101001;
DRAM[57385] = 8'b11101000;
DRAM[57386] = 8'b11100110;
DRAM[57387] = 8'b11100101;
DRAM[57388] = 8'b11100100;
DRAM[57389] = 8'b11100100;
DRAM[57390] = 8'b11100100;
DRAM[57391] = 8'b11100100;
DRAM[57392] = 8'b11011101;
DRAM[57393] = 8'b11100111;
DRAM[57394] = 8'b11100100;
DRAM[57395] = 8'b11010100;
DRAM[57396] = 8'b11001010;
DRAM[57397] = 8'b11001011;
DRAM[57398] = 8'b11000100;
DRAM[57399] = 8'b10110110;
DRAM[57400] = 8'b10110010;
DRAM[57401] = 8'b10101001;
DRAM[57402] = 8'b10100010;
DRAM[57403] = 8'b10100001;
DRAM[57404] = 8'b10100010;
DRAM[57405] = 8'b10100100;
DRAM[57406] = 8'b10101001;
DRAM[57407] = 8'b10101110;
DRAM[57408] = 8'b10101111;
DRAM[57409] = 8'b10110101;
DRAM[57410] = 8'b10111001;
DRAM[57411] = 8'b10110110;
DRAM[57412] = 8'b10101101;
DRAM[57413] = 8'b10100011;
DRAM[57414] = 8'b10011111;
DRAM[57415] = 8'b10011110;
DRAM[57416] = 8'b10010011;
DRAM[57417] = 8'b10011001;
DRAM[57418] = 8'b10100000;
DRAM[57419] = 8'b10100001;
DRAM[57420] = 8'b10011001;
DRAM[57421] = 8'b10010000;
DRAM[57422] = 8'b10010011;
DRAM[57423] = 8'b10011011;
DRAM[57424] = 8'b10011010;
DRAM[57425] = 8'b10100011;
DRAM[57426] = 8'b10000110;
DRAM[57427] = 8'b10001010;
DRAM[57428] = 8'b10001011;
DRAM[57429] = 8'b10010000;
DRAM[57430] = 8'b10000110;
DRAM[57431] = 8'b10100111;
DRAM[57432] = 8'b1111101;
DRAM[57433] = 8'b10011100;
DRAM[57434] = 8'b10010101;
DRAM[57435] = 8'b10000100;
DRAM[57436] = 8'b10010011;
DRAM[57437] = 8'b10010011;
DRAM[57438] = 8'b10000100;
DRAM[57439] = 8'b10001000;
DRAM[57440] = 8'b1111011;
DRAM[57441] = 8'b10000011;
DRAM[57442] = 8'b10001000;
DRAM[57443] = 8'b10000101;
DRAM[57444] = 8'b1111101;
DRAM[57445] = 8'b1111010;
DRAM[57446] = 8'b1111100;
DRAM[57447] = 8'b10000000;
DRAM[57448] = 8'b1101001;
DRAM[57449] = 8'b1110111;
DRAM[57450] = 8'b1101110;
DRAM[57451] = 8'b1100110;
DRAM[57452] = 8'b1110011;
DRAM[57453] = 8'b1110011;
DRAM[57454] = 8'b1100011;
DRAM[57455] = 8'b1100000;
DRAM[57456] = 8'b1101100;
DRAM[57457] = 8'b1100111;
DRAM[57458] = 8'b1101001;
DRAM[57459] = 8'b1100111;
DRAM[57460] = 8'b1100010;
DRAM[57461] = 8'b1100101;
DRAM[57462] = 8'b1100000;
DRAM[57463] = 8'b1001110;
DRAM[57464] = 8'b1100001;
DRAM[57465] = 8'b1100011;
DRAM[57466] = 8'b1100000;
DRAM[57467] = 8'b1011100;
DRAM[57468] = 8'b1100100;
DRAM[57469] = 8'b1110010;
DRAM[57470] = 8'b1110001;
DRAM[57471] = 8'b1100111;
DRAM[57472] = 8'b1101001;
DRAM[57473] = 8'b1101110;
DRAM[57474] = 8'b1110000;
DRAM[57475] = 8'b1101001;
DRAM[57476] = 8'b1100000;
DRAM[57477] = 8'b1011111;
DRAM[57478] = 8'b1100111;
DRAM[57479] = 8'b1110000;
DRAM[57480] = 8'b1011110;
DRAM[57481] = 8'b1011010;
DRAM[57482] = 8'b1011110;
DRAM[57483] = 8'b1101001;
DRAM[57484] = 8'b1101110;
DRAM[57485] = 8'b1101001;
DRAM[57486] = 8'b1100100;
DRAM[57487] = 8'b1100011;
DRAM[57488] = 8'b1101011;
DRAM[57489] = 8'b1100110;
DRAM[57490] = 8'b1101000;
DRAM[57491] = 8'b1110001;
DRAM[57492] = 8'b1110100;
DRAM[57493] = 8'b1101101;
DRAM[57494] = 8'b1101100;
DRAM[57495] = 8'b1110000;
DRAM[57496] = 8'b1100011;
DRAM[57497] = 8'b1101101;
DRAM[57498] = 8'b1110001;
DRAM[57499] = 8'b1101110;
DRAM[57500] = 8'b1110100;
DRAM[57501] = 8'b10000011;
DRAM[57502] = 8'b10001000;
DRAM[57503] = 8'b10000001;
DRAM[57504] = 8'b10001100;
DRAM[57505] = 8'b10010001;
DRAM[57506] = 8'b10010001;
DRAM[57507] = 8'b10001000;
DRAM[57508] = 8'b10000011;
DRAM[57509] = 8'b10001011;
DRAM[57510] = 8'b10011100;
DRAM[57511] = 8'b10100111;
DRAM[57512] = 8'b10010101;
DRAM[57513] = 8'b10011010;
DRAM[57514] = 8'b10011110;
DRAM[57515] = 8'b10011101;
DRAM[57516] = 8'b10100000;
DRAM[57517] = 8'b10100111;
DRAM[57518] = 8'b10101100;
DRAM[57519] = 8'b10101101;
DRAM[57520] = 8'b10101000;
DRAM[57521] = 8'b10101100;
DRAM[57522] = 8'b10110001;
DRAM[57523] = 8'b10110110;
DRAM[57524] = 8'b10111010;
DRAM[57525] = 8'b10111110;
DRAM[57526] = 8'b11000010;
DRAM[57527] = 8'b11000101;
DRAM[57528] = 8'b11010000;
DRAM[57529] = 8'b11010100;
DRAM[57530] = 8'b11011011;
DRAM[57531] = 8'b11100011;
DRAM[57532] = 8'b11101011;
DRAM[57533] = 8'b11110010;
DRAM[57534] = 8'b11110111;
DRAM[57535] = 8'b11111001;
DRAM[57536] = 8'b11111001;
DRAM[57537] = 8'b11111010;
DRAM[57538] = 8'b11100101;
DRAM[57539] = 8'b10111110;
DRAM[57540] = 8'b10100010;
DRAM[57541] = 8'b10011010;
DRAM[57542] = 8'b10010101;
DRAM[57543] = 8'b10001011;
DRAM[57544] = 8'b10001101;
DRAM[57545] = 8'b10000111;
DRAM[57546] = 8'b10000101;
DRAM[57547] = 8'b10000111;
DRAM[57548] = 8'b10000111;
DRAM[57549] = 8'b10000100;
DRAM[57550] = 8'b10000010;
DRAM[57551] = 8'b10000100;
DRAM[57552] = 8'b10000000;
DRAM[57553] = 8'b1111111;
DRAM[57554] = 8'b1111101;
DRAM[57555] = 8'b1111010;
DRAM[57556] = 8'b1111000;
DRAM[57557] = 8'b1110111;
DRAM[57558] = 8'b1110110;
DRAM[57559] = 8'b1110110;
DRAM[57560] = 8'b1110111;
DRAM[57561] = 8'b1110110;
DRAM[57562] = 8'b1110100;
DRAM[57563] = 8'b1110100;
DRAM[57564] = 8'b1110100;
DRAM[57565] = 8'b1110100;
DRAM[57566] = 8'b1110010;
DRAM[57567] = 8'b1110001;
DRAM[57568] = 8'b1101110;
DRAM[57569] = 8'b1101100;
DRAM[57570] = 8'b1101011;
DRAM[57571] = 8'b1101001;
DRAM[57572] = 8'b1101001;
DRAM[57573] = 8'b1101010;
DRAM[57574] = 8'b1101011;
DRAM[57575] = 8'b1101011;
DRAM[57576] = 8'b1101100;
DRAM[57577] = 8'b1101010;
DRAM[57578] = 8'b1101000;
DRAM[57579] = 8'b1101000;
DRAM[57580] = 8'b1101001;
DRAM[57581] = 8'b1101001;
DRAM[57582] = 8'b1101000;
DRAM[57583] = 8'b1100111;
DRAM[57584] = 8'b1101000;
DRAM[57585] = 8'b1101000;
DRAM[57586] = 8'b1101001;
DRAM[57587] = 8'b1101001;
DRAM[57588] = 8'b1101010;
DRAM[57589] = 8'b1101011;
DRAM[57590] = 8'b1101100;
DRAM[57591] = 8'b1101100;
DRAM[57592] = 8'b1101000;
DRAM[57593] = 8'b1101001;
DRAM[57594] = 8'b1101010;
DRAM[57595] = 8'b1101011;
DRAM[57596] = 8'b1101010;
DRAM[57597] = 8'b1101001;
DRAM[57598] = 8'b1101000;
DRAM[57599] = 8'b1100111;
DRAM[57600] = 8'b10001110;
DRAM[57601] = 8'b10001101;
DRAM[57602] = 8'b10001100;
DRAM[57603] = 8'b10001011;
DRAM[57604] = 8'b10001011;
DRAM[57605] = 8'b10001101;
DRAM[57606] = 8'b10010000;
DRAM[57607] = 8'b10010001;
DRAM[57608] = 8'b10010101;
DRAM[57609] = 8'b10010101;
DRAM[57610] = 8'b10011000;
DRAM[57611] = 8'b10011101;
DRAM[57612] = 8'b10011110;
DRAM[57613] = 8'b10100001;
DRAM[57614] = 8'b10101010;
DRAM[57615] = 8'b10110100;
DRAM[57616] = 8'b11001010;
DRAM[57617] = 8'b11100010;
DRAM[57618] = 8'b11110111;
DRAM[57619] = 8'b11111100;
DRAM[57620] = 8'b11111011;
DRAM[57621] = 8'b11111110;
DRAM[57622] = 8'b11111110;
DRAM[57623] = 8'b11111010;
DRAM[57624] = 8'b11111011;
DRAM[57625] = 8'b11111000;
DRAM[57626] = 8'b11110101;
DRAM[57627] = 8'b11110011;
DRAM[57628] = 8'b11110010;
DRAM[57629] = 8'b11110000;
DRAM[57630] = 8'b11101100;
DRAM[57631] = 8'b11101010;
DRAM[57632] = 8'b11110000;
DRAM[57633] = 8'b11110010;
DRAM[57634] = 8'b11110100;
DRAM[57635] = 8'b11110100;
DRAM[57636] = 8'b11110010;
DRAM[57637] = 8'b11101111;
DRAM[57638] = 8'b11101110;
DRAM[57639] = 8'b11101110;
DRAM[57640] = 8'b11101011;
DRAM[57641] = 8'b11101000;
DRAM[57642] = 8'b11100110;
DRAM[57643] = 8'b11100110;
DRAM[57644] = 8'b11100111;
DRAM[57645] = 8'b11100111;
DRAM[57646] = 8'b11100101;
DRAM[57647] = 8'b11100011;
DRAM[57648] = 8'b11011111;
DRAM[57649] = 8'b11010110;
DRAM[57650] = 8'b11010011;
DRAM[57651] = 8'b11010110;
DRAM[57652] = 8'b11010001;
DRAM[57653] = 8'b11000100;
DRAM[57654] = 8'b10111111;
DRAM[57655] = 8'b11000011;
DRAM[57656] = 8'b10110000;
DRAM[57657] = 8'b10110010;
DRAM[57658] = 8'b10110101;
DRAM[57659] = 8'b10110011;
DRAM[57660] = 8'b10101100;
DRAM[57661] = 8'b10101001;
DRAM[57662] = 8'b10110011;
DRAM[57663] = 8'b11000000;
DRAM[57664] = 8'b10110110;
DRAM[57665] = 8'b10111000;
DRAM[57666] = 8'b10111000;
DRAM[57667] = 8'b10110100;
DRAM[57668] = 8'b10101011;
DRAM[57669] = 8'b10100100;
DRAM[57670] = 8'b10100000;
DRAM[57671] = 8'b10011111;
DRAM[57672] = 8'b10011100;
DRAM[57673] = 8'b10011000;
DRAM[57674] = 8'b10010110;
DRAM[57675] = 8'b10010101;
DRAM[57676] = 8'b10010010;
DRAM[57677] = 8'b10010010;
DRAM[57678] = 8'b10011001;
DRAM[57679] = 8'b10100010;
DRAM[57680] = 8'b10011111;
DRAM[57681] = 8'b10001010;
DRAM[57682] = 8'b10001110;
DRAM[57683] = 8'b10011011;
DRAM[57684] = 8'b10000011;
DRAM[57685] = 8'b10001001;
DRAM[57686] = 8'b10010010;
DRAM[57687] = 8'b10001101;
DRAM[57688] = 8'b10000010;
DRAM[57689] = 8'b10010111;
DRAM[57690] = 8'b10001011;
DRAM[57691] = 8'b1111111;
DRAM[57692] = 8'b10010000;
DRAM[57693] = 8'b10001111;
DRAM[57694] = 8'b10000001;
DRAM[57695] = 8'b10000111;
DRAM[57696] = 8'b10000010;
DRAM[57697] = 8'b10000110;
DRAM[57698] = 8'b10000101;
DRAM[57699] = 8'b10000000;
DRAM[57700] = 8'b1111110;
DRAM[57701] = 8'b10000000;
DRAM[57702] = 8'b1111111;
DRAM[57703] = 8'b1111011;
DRAM[57704] = 8'b1101110;
DRAM[57705] = 8'b1110001;
DRAM[57706] = 8'b1101011;
DRAM[57707] = 8'b1101010;
DRAM[57708] = 8'b1110011;
DRAM[57709] = 8'b1110100;
DRAM[57710] = 8'b1101010;
DRAM[57711] = 8'b1100101;
DRAM[57712] = 8'b1101110;
DRAM[57713] = 8'b1101001;
DRAM[57714] = 8'b1101001;
DRAM[57715] = 8'b1100101;
DRAM[57716] = 8'b1011111;
DRAM[57717] = 8'b1100100;
DRAM[57718] = 8'b1100100;
DRAM[57719] = 8'b1010111;
DRAM[57720] = 8'b1100011;
DRAM[57721] = 8'b1100111;
DRAM[57722] = 8'b1100111;
DRAM[57723] = 8'b1100100;
DRAM[57724] = 8'b1101010;
DRAM[57725] = 8'b1110011;
DRAM[57726] = 8'b1110010;
DRAM[57727] = 8'b1101000;
DRAM[57728] = 8'b1100110;
DRAM[57729] = 8'b1110000;
DRAM[57730] = 8'b1110100;
DRAM[57731] = 8'b1101100;
DRAM[57732] = 8'b1100011;
DRAM[57733] = 8'b1100100;
DRAM[57734] = 8'b1101010;
DRAM[57735] = 8'b1101101;
DRAM[57736] = 8'b1101010;
DRAM[57737] = 8'b1100001;
DRAM[57738] = 8'b1011101;
DRAM[57739] = 8'b1100110;
DRAM[57740] = 8'b1101111;
DRAM[57741] = 8'b1101111;
DRAM[57742] = 8'b1101011;
DRAM[57743] = 8'b1101000;
DRAM[57744] = 8'b1100111;
DRAM[57745] = 8'b1100110;
DRAM[57746] = 8'b1101000;
DRAM[57747] = 8'b1101111;
DRAM[57748] = 8'b1110010;
DRAM[57749] = 8'b1110001;
DRAM[57750] = 8'b1110001;
DRAM[57751] = 8'b1110011;
DRAM[57752] = 8'b1111000;
DRAM[57753] = 8'b1101111;
DRAM[57754] = 8'b1101111;
DRAM[57755] = 8'b1111000;
DRAM[57756] = 8'b1111011;
DRAM[57757] = 8'b1110101;
DRAM[57758] = 8'b1110111;
DRAM[57759] = 8'b10000000;
DRAM[57760] = 8'b1111110;
DRAM[57761] = 8'b10000110;
DRAM[57762] = 8'b10001011;
DRAM[57763] = 8'b10001100;
DRAM[57764] = 8'b10001100;
DRAM[57765] = 8'b10001111;
DRAM[57766] = 8'b10001111;
DRAM[57767] = 8'b10001101;
DRAM[57768] = 8'b10010111;
DRAM[57769] = 8'b10011011;
DRAM[57770] = 8'b10011011;
DRAM[57771] = 8'b10011001;
DRAM[57772] = 8'b10011100;
DRAM[57773] = 8'b10100101;
DRAM[57774] = 8'b10101101;
DRAM[57775] = 8'b10110000;
DRAM[57776] = 8'b10101110;
DRAM[57777] = 8'b10110001;
DRAM[57778] = 8'b10110101;
DRAM[57779] = 8'b10111000;
DRAM[57780] = 8'b10111011;
DRAM[57781] = 8'b10111110;
DRAM[57782] = 8'b11000010;
DRAM[57783] = 8'b11000101;
DRAM[57784] = 8'b11010100;
DRAM[57785] = 8'b11010111;
DRAM[57786] = 8'b11011101;
DRAM[57787] = 8'b11100101;
DRAM[57788] = 8'b11101101;
DRAM[57789] = 8'b11110101;
DRAM[57790] = 8'b11111010;
DRAM[57791] = 8'b11111101;
DRAM[57792] = 8'b11110111;
DRAM[57793] = 8'b11111010;
DRAM[57794] = 8'b11101001;
DRAM[57795] = 8'b11000101;
DRAM[57796] = 8'b10101001;
DRAM[57797] = 8'b10011110;
DRAM[57798] = 8'b10010101;
DRAM[57799] = 8'b10001010;
DRAM[57800] = 8'b10001100;
DRAM[57801] = 8'b10000111;
DRAM[57802] = 8'b10000100;
DRAM[57803] = 8'b10000110;
DRAM[57804] = 8'b10000111;
DRAM[57805] = 8'b10000100;
DRAM[57806] = 8'b10000011;
DRAM[57807] = 8'b10000100;
DRAM[57808] = 8'b10000001;
DRAM[57809] = 8'b10000000;
DRAM[57810] = 8'b1111101;
DRAM[57811] = 8'b1111011;
DRAM[57812] = 8'b1111001;
DRAM[57813] = 8'b1111000;
DRAM[57814] = 8'b1110111;
DRAM[57815] = 8'b1110110;
DRAM[57816] = 8'b1110111;
DRAM[57817] = 8'b1110101;
DRAM[57818] = 8'b1110011;
DRAM[57819] = 8'b1110100;
DRAM[57820] = 8'b1110100;
DRAM[57821] = 8'b1110101;
DRAM[57822] = 8'b1110011;
DRAM[57823] = 8'b1110001;
DRAM[57824] = 8'b1101110;
DRAM[57825] = 8'b1101101;
DRAM[57826] = 8'b1101011;
DRAM[57827] = 8'b1101010;
DRAM[57828] = 8'b1101010;
DRAM[57829] = 8'b1101010;
DRAM[57830] = 8'b1101011;
DRAM[57831] = 8'b1101100;
DRAM[57832] = 8'b1101100;
DRAM[57833] = 8'b1101010;
DRAM[57834] = 8'b1101000;
DRAM[57835] = 8'b1101000;
DRAM[57836] = 8'b1101001;
DRAM[57837] = 8'b1101001;
DRAM[57838] = 8'b1101001;
DRAM[57839] = 8'b1100111;
DRAM[57840] = 8'b1101000;
DRAM[57841] = 8'b1101000;
DRAM[57842] = 8'b1101001;
DRAM[57843] = 8'b1101010;
DRAM[57844] = 8'b1101011;
DRAM[57845] = 8'b1101011;
DRAM[57846] = 8'b1101100;
DRAM[57847] = 8'b1101100;
DRAM[57848] = 8'b1101001;
DRAM[57849] = 8'b1101010;
DRAM[57850] = 8'b1101011;
DRAM[57851] = 8'b1101011;
DRAM[57852] = 8'b1101011;
DRAM[57853] = 8'b1101010;
DRAM[57854] = 8'b1101000;
DRAM[57855] = 8'b1100111;
DRAM[57856] = 8'b10001010;
DRAM[57857] = 8'b10001010;
DRAM[57858] = 8'b10001010;
DRAM[57859] = 8'b10001011;
DRAM[57860] = 8'b10001100;
DRAM[57861] = 8'b10001101;
DRAM[57862] = 8'b10001111;
DRAM[57863] = 8'b10010000;
DRAM[57864] = 8'b10010011;
DRAM[57865] = 8'b10010101;
DRAM[57866] = 8'b10011001;
DRAM[57867] = 8'b10011100;
DRAM[57868] = 8'b10011100;
DRAM[57869] = 8'b10011111;
DRAM[57870] = 8'b10101100;
DRAM[57871] = 8'b10111010;
DRAM[57872] = 8'b11011000;
DRAM[57873] = 8'b11101011;
DRAM[57874] = 8'b11111100;
DRAM[57875] = 8'b11111111;
DRAM[57876] = 8'b11111110;
DRAM[57877] = 8'b11111111;
DRAM[57878] = 8'b11111110;
DRAM[57879] = 8'b11111010;
DRAM[57880] = 8'b11111001;
DRAM[57881] = 8'b11110111;
DRAM[57882] = 8'b11110101;
DRAM[57883] = 8'b11110011;
DRAM[57884] = 8'b11110001;
DRAM[57885] = 8'b11101101;
DRAM[57886] = 8'b11101000;
DRAM[57887] = 8'b11100100;
DRAM[57888] = 8'b11101111;
DRAM[57889] = 8'b11101110;
DRAM[57890] = 8'b11101110;
DRAM[57891] = 8'b11101111;
DRAM[57892] = 8'b11110000;
DRAM[57893] = 8'b11101110;
DRAM[57894] = 8'b11101100;
DRAM[57895] = 8'b11101001;
DRAM[57896] = 8'b11101000;
DRAM[57897] = 8'b11100100;
DRAM[57898] = 8'b11100001;
DRAM[57899] = 8'b11100010;
DRAM[57900] = 8'b11100110;
DRAM[57901] = 8'b11100111;
DRAM[57902] = 8'b11100010;
DRAM[57903] = 8'b11011110;
DRAM[57904] = 8'b11011001;
DRAM[57905] = 8'b11001100;
DRAM[57906] = 8'b11000111;
DRAM[57907] = 8'b11001110;
DRAM[57908] = 8'b11001101;
DRAM[57909] = 8'b11000010;
DRAM[57910] = 8'b10111101;
DRAM[57911] = 8'b11000010;
DRAM[57912] = 8'b10110010;
DRAM[57913] = 8'b10101011;
DRAM[57914] = 8'b10101010;
DRAM[57915] = 8'b10110011;
DRAM[57916] = 8'b10111101;
DRAM[57917] = 8'b11000000;
DRAM[57918] = 8'b10111110;
DRAM[57919] = 8'b10111101;
DRAM[57920] = 8'b10110101;
DRAM[57921] = 8'b10110100;
DRAM[57922] = 8'b10110011;
DRAM[57923] = 8'b10110001;
DRAM[57924] = 8'b10101111;
DRAM[57925] = 8'b10101101;
DRAM[57926] = 8'b10101100;
DRAM[57927] = 8'b10101011;
DRAM[57928] = 8'b10100101;
DRAM[57929] = 8'b10011100;
DRAM[57930] = 8'b10010101;
DRAM[57931] = 8'b10010010;
DRAM[57932] = 8'b10010001;
DRAM[57933] = 8'b10010000;
DRAM[57934] = 8'b10010100;
DRAM[57935] = 8'b10011001;
DRAM[57936] = 8'b10011100;
DRAM[57937] = 8'b10000010;
DRAM[57938] = 8'b10001110;
DRAM[57939] = 8'b10010011;
DRAM[57940] = 8'b10000111;
DRAM[57941] = 8'b10000001;
DRAM[57942] = 8'b10001110;
DRAM[57943] = 8'b10000001;
DRAM[57944] = 8'b10001100;
DRAM[57945] = 8'b10010010;
DRAM[57946] = 8'b10000100;
DRAM[57947] = 8'b1111111;
DRAM[57948] = 8'b10001110;
DRAM[57949] = 8'b10001010;
DRAM[57950] = 8'b1111111;
DRAM[57951] = 8'b10000111;
DRAM[57952] = 8'b10001010;
DRAM[57953] = 8'b10001011;
DRAM[57954] = 8'b10000100;
DRAM[57955] = 8'b1111010;
DRAM[57956] = 8'b1111101;
DRAM[57957] = 8'b10000110;
DRAM[57958] = 8'b10000010;
DRAM[57959] = 8'b1110110;
DRAM[57960] = 8'b1111011;
DRAM[57961] = 8'b1101101;
DRAM[57962] = 8'b1101011;
DRAM[57963] = 8'b1110001;
DRAM[57964] = 8'b1110011;
DRAM[57965] = 8'b1110100;
DRAM[57966] = 8'b1110001;
DRAM[57967] = 8'b1101000;
DRAM[57968] = 8'b1110000;
DRAM[57969] = 8'b1101010;
DRAM[57970] = 8'b1101001;
DRAM[57971] = 8'b1100101;
DRAM[57972] = 8'b1011101;
DRAM[57973] = 8'b1100011;
DRAM[57974] = 8'b1101001;
DRAM[57975] = 8'b1100010;
DRAM[57976] = 8'b1100011;
DRAM[57977] = 8'b1101010;
DRAM[57978] = 8'b1101110;
DRAM[57979] = 8'b1101011;
DRAM[57980] = 8'b1101100;
DRAM[57981] = 8'b1110001;
DRAM[57982] = 8'b1101111;
DRAM[57983] = 8'b1101000;
DRAM[57984] = 8'b1100011;
DRAM[57985] = 8'b1110011;
DRAM[57986] = 8'b1111001;
DRAM[57987] = 8'b1101101;
DRAM[57988] = 8'b1100100;
DRAM[57989] = 8'b1101001;
DRAM[57990] = 8'b1101101;
DRAM[57991] = 8'b1101011;
DRAM[57992] = 8'b1110100;
DRAM[57993] = 8'b1100110;
DRAM[57994] = 8'b1011100;
DRAM[57995] = 8'b1100001;
DRAM[57996] = 8'b1101101;
DRAM[57997] = 8'b1110010;
DRAM[57998] = 8'b1110000;
DRAM[57999] = 8'b1101100;
DRAM[58000] = 8'b1100101;
DRAM[58001] = 8'b1101001;
DRAM[58002] = 8'b1101100;
DRAM[58003] = 8'b1101100;
DRAM[58004] = 8'b1101111;
DRAM[58005] = 8'b1110100;
DRAM[58006] = 8'b1110101;
DRAM[58007] = 8'b1110011;
DRAM[58008] = 8'b1111110;
DRAM[58009] = 8'b1110011;
DRAM[58010] = 8'b1110001;
DRAM[58011] = 8'b1111010;
DRAM[58012] = 8'b1111100;
DRAM[58013] = 8'b1110110;
DRAM[58014] = 8'b1110110;
DRAM[58015] = 8'b1111110;
DRAM[58016] = 8'b1111001;
DRAM[58017] = 8'b1111110;
DRAM[58018] = 8'b10000100;
DRAM[58019] = 8'b10001010;
DRAM[58020] = 8'b10010001;
DRAM[58021] = 8'b10010011;
DRAM[58022] = 8'b10001100;
DRAM[58023] = 8'b10000010;
DRAM[58024] = 8'b10001100;
DRAM[58025] = 8'b10010100;
DRAM[58026] = 8'b10011011;
DRAM[58027] = 8'b10011101;
DRAM[58028] = 8'b10100000;
DRAM[58029] = 8'b10100100;
DRAM[58030] = 8'b10100101;
DRAM[58031] = 8'b10100011;
DRAM[58032] = 8'b10101000;
DRAM[58033] = 8'b10101010;
DRAM[58034] = 8'b10101101;
DRAM[58035] = 8'b10110000;
DRAM[58036] = 8'b10110011;
DRAM[58037] = 8'b10110111;
DRAM[58038] = 8'b10111101;
DRAM[58039] = 8'b11000001;
DRAM[58040] = 8'b11001111;
DRAM[58041] = 8'b11010011;
DRAM[58042] = 8'b11011010;
DRAM[58043] = 8'b11100011;
DRAM[58044] = 8'b11101011;
DRAM[58045] = 8'b11110010;
DRAM[58046] = 8'b11110111;
DRAM[58047] = 8'b11111001;
DRAM[58048] = 8'b11110101;
DRAM[58049] = 8'b11110111;
DRAM[58050] = 8'b11101001;
DRAM[58051] = 8'b11001000;
DRAM[58052] = 8'b10101100;
DRAM[58053] = 8'b10011111;
DRAM[58054] = 8'b10010011;
DRAM[58055] = 8'b10001000;
DRAM[58056] = 8'b10001011;
DRAM[58057] = 8'b10000110;
DRAM[58058] = 8'b10000011;
DRAM[58059] = 8'b10000110;
DRAM[58060] = 8'b10000111;
DRAM[58061] = 8'b10000100;
DRAM[58062] = 8'b10000011;
DRAM[58063] = 8'b10000101;
DRAM[58064] = 8'b10000001;
DRAM[58065] = 8'b10000000;
DRAM[58066] = 8'b1111110;
DRAM[58067] = 8'b1111011;
DRAM[58068] = 8'b1111001;
DRAM[58069] = 8'b1111000;
DRAM[58070] = 8'b1110111;
DRAM[58071] = 8'b1110111;
DRAM[58072] = 8'b1110110;
DRAM[58073] = 8'b1110100;
DRAM[58074] = 8'b1110011;
DRAM[58075] = 8'b1110011;
DRAM[58076] = 8'b1110101;
DRAM[58077] = 8'b1110101;
DRAM[58078] = 8'b1110100;
DRAM[58079] = 8'b1110010;
DRAM[58080] = 8'b1101111;
DRAM[58081] = 8'b1101110;
DRAM[58082] = 8'b1101100;
DRAM[58083] = 8'b1101011;
DRAM[58084] = 8'b1101010;
DRAM[58085] = 8'b1101011;
DRAM[58086] = 8'b1101100;
DRAM[58087] = 8'b1101101;
DRAM[58088] = 8'b1101100;
DRAM[58089] = 8'b1101010;
DRAM[58090] = 8'b1101000;
DRAM[58091] = 8'b1101000;
DRAM[58092] = 8'b1101001;
DRAM[58093] = 8'b1101010;
DRAM[58094] = 8'b1101001;
DRAM[58095] = 8'b1101000;
DRAM[58096] = 8'b1101001;
DRAM[58097] = 8'b1101001;
DRAM[58098] = 8'b1101010;
DRAM[58099] = 8'b1101010;
DRAM[58100] = 8'b1101011;
DRAM[58101] = 8'b1101100;
DRAM[58102] = 8'b1101101;
DRAM[58103] = 8'b1101101;
DRAM[58104] = 8'b1101011;
DRAM[58105] = 8'b1101100;
DRAM[58106] = 8'b1101100;
DRAM[58107] = 8'b1101100;
DRAM[58108] = 8'b1101100;
DRAM[58109] = 8'b1101011;
DRAM[58110] = 8'b1101001;
DRAM[58111] = 8'b1101001;
DRAM[58112] = 8'b10000111;
DRAM[58113] = 8'b10001000;
DRAM[58114] = 8'b10001001;
DRAM[58115] = 8'b10001010;
DRAM[58116] = 8'b10001100;
DRAM[58117] = 8'b10001101;
DRAM[58118] = 8'b10001110;
DRAM[58119] = 8'b10001111;
DRAM[58120] = 8'b10010011;
DRAM[58121] = 8'b10010101;
DRAM[58122] = 8'b10011000;
DRAM[58123] = 8'b10011001;
DRAM[58124] = 8'b10010111;
DRAM[58125] = 8'b10011010;
DRAM[58126] = 8'b10101010;
DRAM[58127] = 8'b10111011;
DRAM[58128] = 8'b11011101;
DRAM[58129] = 8'b11101100;
DRAM[58130] = 8'b11111001;
DRAM[58131] = 8'b11111101;
DRAM[58132] = 8'b11111110;
DRAM[58133] = 8'b11111111;
DRAM[58134] = 8'b11111110;
DRAM[58135] = 8'b11111011;
DRAM[58136] = 8'b11111011;
DRAM[58137] = 8'b11111000;
DRAM[58138] = 8'b11110100;
DRAM[58139] = 8'b11110010;
DRAM[58140] = 8'b11110000;
DRAM[58141] = 8'b11101101;
DRAM[58142] = 8'b11101010;
DRAM[58143] = 8'b11100111;
DRAM[58144] = 8'b11101100;
DRAM[58145] = 8'b11101010;
DRAM[58146] = 8'b11101001;
DRAM[58147] = 8'b11101011;
DRAM[58148] = 8'b11101110;
DRAM[58149] = 8'b11101110;
DRAM[58150] = 8'b11101010;
DRAM[58151] = 8'b11100110;
DRAM[58152] = 8'b11100001;
DRAM[58153] = 8'b11011100;
DRAM[58154] = 8'b11011000;
DRAM[58155] = 8'b11011011;
DRAM[58156] = 8'b11100000;
DRAM[58157] = 8'b11100000;
DRAM[58158] = 8'b11011001;
DRAM[58159] = 8'b11010010;
DRAM[58160] = 8'b11001011;
DRAM[58161] = 8'b11001101;
DRAM[58162] = 8'b11001001;
DRAM[58163] = 8'b11000010;
DRAM[58164] = 8'b11000011;
DRAM[58165] = 8'b11001000;
DRAM[58166] = 8'b11000001;
DRAM[58167] = 8'b10110101;
DRAM[58168] = 8'b10111001;
DRAM[58169] = 8'b10110000;
DRAM[58170] = 8'b10101110;
DRAM[58171] = 8'b10111000;
DRAM[58172] = 8'b11000011;
DRAM[58173] = 8'b11000011;
DRAM[58174] = 8'b10111010;
DRAM[58175] = 8'b10110010;
DRAM[58176] = 8'b10110010;
DRAM[58177] = 8'b10110000;
DRAM[58178] = 8'b10101110;
DRAM[58179] = 8'b10101101;
DRAM[58180] = 8'b10101100;
DRAM[58181] = 8'b10101010;
DRAM[58182] = 8'b10100111;
DRAM[58183] = 8'b10100101;
DRAM[58184] = 8'b10011001;
DRAM[58185] = 8'b10010110;
DRAM[58186] = 8'b10010101;
DRAM[58187] = 8'b10010111;
DRAM[58188] = 8'b10010101;
DRAM[58189] = 8'b10010000;
DRAM[58190] = 8'b10001101;
DRAM[58191] = 8'b10001110;
DRAM[58192] = 8'b10010000;
DRAM[58193] = 8'b10001111;
DRAM[58194] = 8'b10000110;
DRAM[58195] = 8'b1110111;
DRAM[58196] = 8'b10010011;
DRAM[58197] = 8'b1111101;
DRAM[58198] = 8'b1111010;
DRAM[58199] = 8'b10001010;
DRAM[58200] = 8'b10001110;
DRAM[58201] = 8'b10001110;
DRAM[58202] = 8'b10000101;
DRAM[58203] = 8'b10000101;
DRAM[58204] = 8'b10001101;
DRAM[58205] = 8'b10000101;
DRAM[58206] = 8'b1111110;
DRAM[58207] = 8'b10001011;
DRAM[58208] = 8'b10001100;
DRAM[58209] = 8'b10001110;
DRAM[58210] = 8'b10000101;
DRAM[58211] = 8'b1111000;
DRAM[58212] = 8'b1111010;
DRAM[58213] = 8'b10000110;
DRAM[58214] = 8'b10000011;
DRAM[58215] = 8'b1110101;
DRAM[58216] = 8'b10001010;
DRAM[58217] = 8'b1101111;
DRAM[58218] = 8'b1101101;
DRAM[58219] = 8'b1111000;
DRAM[58220] = 8'b1110010;
DRAM[58221] = 8'b1110010;
DRAM[58222] = 8'b1110011;
DRAM[58223] = 8'b1101000;
DRAM[58224] = 8'b1101110;
DRAM[58225] = 8'b1101000;
DRAM[58226] = 8'b1101001;
DRAM[58227] = 8'b1100110;
DRAM[58228] = 8'b1011110;
DRAM[58229] = 8'b1100011;
DRAM[58230] = 8'b1101011;
DRAM[58231] = 8'b1101001;
DRAM[58232] = 8'b1100011;
DRAM[58233] = 8'b1101011;
DRAM[58234] = 8'b1101111;
DRAM[58235] = 8'b1101100;
DRAM[58236] = 8'b1101010;
DRAM[58237] = 8'b1101011;
DRAM[58238] = 8'b1101011;
DRAM[58239] = 8'b1101000;
DRAM[58240] = 8'b1100011;
DRAM[58241] = 8'b1110100;
DRAM[58242] = 8'b1111001;
DRAM[58243] = 8'b1101011;
DRAM[58244] = 8'b1100011;
DRAM[58245] = 8'b1101010;
DRAM[58246] = 8'b1101111;
DRAM[58247] = 8'b1101100;
DRAM[58248] = 8'b1110011;
DRAM[58249] = 8'b1100111;
DRAM[58250] = 8'b1011101;
DRAM[58251] = 8'b1011110;
DRAM[58252] = 8'b1101000;
DRAM[58253] = 8'b1101111;
DRAM[58254] = 8'b1101111;
DRAM[58255] = 8'b1101100;
DRAM[58256] = 8'b1100110;
DRAM[58257] = 8'b1101110;
DRAM[58258] = 8'b1110000;
DRAM[58259] = 8'b1101011;
DRAM[58260] = 8'b1101100;
DRAM[58261] = 8'b1110101;
DRAM[58262] = 8'b1110111;
DRAM[58263] = 8'b1110011;
DRAM[58264] = 8'b1110001;
DRAM[58265] = 8'b1110111;
DRAM[58266] = 8'b1110111;
DRAM[58267] = 8'b1110001;
DRAM[58268] = 8'b1110111;
DRAM[58269] = 8'b10000100;
DRAM[58270] = 8'b10000110;
DRAM[58271] = 8'b1111101;
DRAM[58272] = 8'b10000001;
DRAM[58273] = 8'b10000001;
DRAM[58274] = 8'b10000000;
DRAM[58275] = 8'b10000001;
DRAM[58276] = 8'b10001000;
DRAM[58277] = 8'b10010001;
DRAM[58278] = 8'b10010011;
DRAM[58279] = 8'b10001111;
DRAM[58280] = 8'b10001011;
DRAM[58281] = 8'b10010010;
DRAM[58282] = 8'b10010111;
DRAM[58283] = 8'b10010111;
DRAM[58284] = 8'b10011001;
DRAM[58285] = 8'b10011101;
DRAM[58286] = 8'b10011110;
DRAM[58287] = 8'b10011101;
DRAM[58288] = 8'b10011110;
DRAM[58289] = 8'b10100001;
DRAM[58290] = 8'b10100100;
DRAM[58291] = 8'b10101000;
DRAM[58292] = 8'b10101101;
DRAM[58293] = 8'b10110100;
DRAM[58294] = 8'b10111011;
DRAM[58295] = 8'b11000001;
DRAM[58296] = 8'b11001010;
DRAM[58297] = 8'b11010000;
DRAM[58298] = 8'b11011001;
DRAM[58299] = 8'b11100100;
DRAM[58300] = 8'b11101100;
DRAM[58301] = 8'b11110010;
DRAM[58302] = 8'b11110100;
DRAM[58303] = 8'b11110101;
DRAM[58304] = 8'b11110101;
DRAM[58305] = 8'b11110100;
DRAM[58306] = 8'b11100011;
DRAM[58307] = 8'b11000010;
DRAM[58308] = 8'b10100110;
DRAM[58309] = 8'b10011001;
DRAM[58310] = 8'b10010001;
DRAM[58311] = 8'b10001001;
DRAM[58312] = 8'b10001011;
DRAM[58313] = 8'b10000110;
DRAM[58314] = 8'b10000100;
DRAM[58315] = 8'b10000110;
DRAM[58316] = 8'b10000111;
DRAM[58317] = 8'b10000101;
DRAM[58318] = 8'b10000100;
DRAM[58319] = 8'b10000110;
DRAM[58320] = 8'b10000000;
DRAM[58321] = 8'b1111111;
DRAM[58322] = 8'b1111101;
DRAM[58323] = 8'b1111011;
DRAM[58324] = 8'b1111000;
DRAM[58325] = 8'b1110111;
DRAM[58326] = 8'b1110110;
DRAM[58327] = 8'b1110110;
DRAM[58328] = 8'b1110101;
DRAM[58329] = 8'b1110100;
DRAM[58330] = 8'b1110011;
DRAM[58331] = 8'b1110011;
DRAM[58332] = 8'b1110101;
DRAM[58333] = 8'b1110101;
DRAM[58334] = 8'b1110100;
DRAM[58335] = 8'b1110011;
DRAM[58336] = 8'b1101111;
DRAM[58337] = 8'b1101110;
DRAM[58338] = 8'b1101100;
DRAM[58339] = 8'b1101011;
DRAM[58340] = 8'b1101011;
DRAM[58341] = 8'b1101011;
DRAM[58342] = 8'b1101100;
DRAM[58343] = 8'b1101101;
DRAM[58344] = 8'b1101011;
DRAM[58345] = 8'b1101001;
DRAM[58346] = 8'b1100111;
DRAM[58347] = 8'b1100111;
DRAM[58348] = 8'b1101001;
DRAM[58349] = 8'b1101010;
DRAM[58350] = 8'b1101001;
DRAM[58351] = 8'b1101000;
DRAM[58352] = 8'b1101010;
DRAM[58353] = 8'b1101010;
DRAM[58354] = 8'b1101010;
DRAM[58355] = 8'b1101011;
DRAM[58356] = 8'b1101100;
DRAM[58357] = 8'b1101101;
DRAM[58358] = 8'b1101101;
DRAM[58359] = 8'b1101110;
DRAM[58360] = 8'b1101101;
DRAM[58361] = 8'b1101101;
DRAM[58362] = 8'b1101101;
DRAM[58363] = 8'b1101101;
DRAM[58364] = 8'b1101100;
DRAM[58365] = 8'b1101011;
DRAM[58366] = 8'b1101010;
DRAM[58367] = 8'b1101010;
DRAM[58368] = 8'b10000111;
DRAM[58369] = 8'b10000111;
DRAM[58370] = 8'b10001001;
DRAM[58371] = 8'b10001010;
DRAM[58372] = 8'b10001011;
DRAM[58373] = 8'b10001101;
DRAM[58374] = 8'b10001110;
DRAM[58375] = 8'b10001110;
DRAM[58376] = 8'b10010011;
DRAM[58377] = 8'b10010100;
DRAM[58378] = 8'b10010111;
DRAM[58379] = 8'b10011000;
DRAM[58380] = 8'b10011000;
DRAM[58381] = 8'b10011111;
DRAM[58382] = 8'b10110011;
DRAM[58383] = 8'b11000110;
DRAM[58384] = 8'b11100101;
DRAM[58385] = 8'b11101110;
DRAM[58386] = 8'b11110111;
DRAM[58387] = 8'b11111100;
DRAM[58388] = 8'b11111101;
DRAM[58389] = 8'b11111111;
DRAM[58390] = 8'b11111110;
DRAM[58391] = 8'b11111100;
DRAM[58392] = 8'b11111101;
DRAM[58393] = 8'b11111000;
DRAM[58394] = 8'b11110011;
DRAM[58395] = 8'b11110000;
DRAM[58396] = 8'b11110000;
DRAM[58397] = 8'b11110000;
DRAM[58398] = 8'b11110001;
DRAM[58399] = 8'b11110000;
DRAM[58400] = 8'b11110010;
DRAM[58401] = 8'b11101111;
DRAM[58402] = 8'b11101101;
DRAM[58403] = 8'b11101101;
DRAM[58404] = 8'b11101110;
DRAM[58405] = 8'b11101100;
DRAM[58406] = 8'b11100111;
DRAM[58407] = 8'b11100010;
DRAM[58408] = 8'b11011010;
DRAM[58409] = 8'b11010110;
DRAM[58410] = 8'b11010011;
DRAM[58411] = 8'b11010101;
DRAM[58412] = 8'b11011010;
DRAM[58413] = 8'b11011001;
DRAM[58414] = 8'b11010000;
DRAM[58415] = 8'b11001000;
DRAM[58416] = 8'b11000100;
DRAM[58417] = 8'b11000110;
DRAM[58418] = 8'b11000101;
DRAM[58419] = 8'b11000011;
DRAM[58420] = 8'b11000111;
DRAM[58421] = 8'b11001010;
DRAM[58422] = 8'b11000011;
DRAM[58423] = 8'b10110111;
DRAM[58424] = 8'b11000011;
DRAM[58425] = 8'b11001010;
DRAM[58426] = 8'b11010000;
DRAM[58427] = 8'b11001101;
DRAM[58428] = 8'b10111110;
DRAM[58429] = 8'b10110000;
DRAM[58430] = 8'b10101111;
DRAM[58431] = 8'b10110110;
DRAM[58432] = 8'b10110101;
DRAM[58433] = 8'b10110011;
DRAM[58434] = 8'b10101110;
DRAM[58435] = 8'b10101001;
DRAM[58436] = 8'b10100011;
DRAM[58437] = 8'b10011011;
DRAM[58438] = 8'b10010010;
DRAM[58439] = 8'b10001101;
DRAM[58440] = 8'b10000111;
DRAM[58441] = 8'b10001001;
DRAM[58442] = 8'b10001111;
DRAM[58443] = 8'b10010011;
DRAM[58444] = 8'b10010000;
DRAM[58445] = 8'b10001010;
DRAM[58446] = 8'b10001001;
DRAM[58447] = 8'b10001110;
DRAM[58448] = 8'b10000111;
DRAM[58449] = 8'b10001000;
DRAM[58450] = 8'b10000011;
DRAM[58451] = 8'b1110110;
DRAM[58452] = 8'b10010011;
DRAM[58453] = 8'b1111100;
DRAM[58454] = 8'b1111010;
DRAM[58455] = 8'b10001010;
DRAM[58456] = 8'b10000010;
DRAM[58457] = 8'b10000010;
DRAM[58458] = 8'b10000100;
DRAM[58459] = 8'b10001001;
DRAM[58460] = 8'b10001010;
DRAM[58461] = 8'b10000001;
DRAM[58462] = 8'b10000011;
DRAM[58463] = 8'b10010010;
DRAM[58464] = 8'b10000111;
DRAM[58465] = 8'b10001100;
DRAM[58466] = 8'b10000111;
DRAM[58467] = 8'b1111010;
DRAM[58468] = 8'b1111000;
DRAM[58469] = 8'b10000000;
DRAM[58470] = 8'b10000000;
DRAM[58471] = 8'b1111000;
DRAM[58472] = 8'b10001101;
DRAM[58473] = 8'b1110010;
DRAM[58474] = 8'b1110000;
DRAM[58475] = 8'b1111010;
DRAM[58476] = 8'b1110100;
DRAM[58477] = 8'b1110100;
DRAM[58478] = 8'b1110111;
DRAM[58479] = 8'b1101110;
DRAM[58480] = 8'b1101011;
DRAM[58481] = 8'b1100101;
DRAM[58482] = 8'b1101001;
DRAM[58483] = 8'b1101010;
DRAM[58484] = 8'b1100011;
DRAM[58485] = 8'b1100101;
DRAM[58486] = 8'b1101101;
DRAM[58487] = 8'b1101011;
DRAM[58488] = 8'b1101000;
DRAM[58489] = 8'b1101110;
DRAM[58490] = 8'b1110001;
DRAM[58491] = 8'b1101101;
DRAM[58492] = 8'b1101001;
DRAM[58493] = 8'b1101001;
DRAM[58494] = 8'b1101010;
DRAM[58495] = 8'b1101011;
DRAM[58496] = 8'b1100101;
DRAM[58497] = 8'b1110011;
DRAM[58498] = 8'b1110110;
DRAM[58499] = 8'b1101000;
DRAM[58500] = 8'b1100000;
DRAM[58501] = 8'b1100111;
DRAM[58502] = 8'b1101111;
DRAM[58503] = 8'b1110000;
DRAM[58504] = 8'b1101110;
DRAM[58505] = 8'b1101001;
DRAM[58506] = 8'b1100011;
DRAM[58507] = 8'b1100010;
DRAM[58508] = 8'b1100111;
DRAM[58509] = 8'b1101100;
DRAM[58510] = 8'b1101101;
DRAM[58511] = 8'b1101011;
DRAM[58512] = 8'b1100110;
DRAM[58513] = 8'b1101111;
DRAM[58514] = 8'b1110001;
DRAM[58515] = 8'b1101011;
DRAM[58516] = 8'b1101100;
DRAM[58517] = 8'b1110110;
DRAM[58518] = 8'b1111010;
DRAM[58519] = 8'b1111000;
DRAM[58520] = 8'b1110001;
DRAM[58521] = 8'b1110111;
DRAM[58522] = 8'b1110111;
DRAM[58523] = 8'b1110011;
DRAM[58524] = 8'b1111010;
DRAM[58525] = 8'b10000111;
DRAM[58526] = 8'b10000110;
DRAM[58527] = 8'b1111100;
DRAM[58528] = 8'b10000101;
DRAM[58529] = 8'b10000100;
DRAM[58530] = 8'b1111111;
DRAM[58531] = 8'b1111000;
DRAM[58532] = 8'b1111010;
DRAM[58533] = 8'b10000101;
DRAM[58534] = 8'b10001111;
DRAM[58535] = 8'b10010100;
DRAM[58536] = 8'b10010110;
DRAM[58537] = 8'b10010111;
DRAM[58538] = 8'b10010011;
DRAM[58539] = 8'b10001100;
DRAM[58540] = 8'b10001101;
DRAM[58541] = 8'b10010110;
DRAM[58542] = 8'b10011111;
DRAM[58543] = 8'b10100011;
DRAM[58544] = 8'b10100001;
DRAM[58545] = 8'b10100011;
DRAM[58546] = 8'b10100111;
DRAM[58547] = 8'b10101011;
DRAM[58548] = 8'b10110000;
DRAM[58549] = 8'b10110111;
DRAM[58550] = 8'b10111111;
DRAM[58551] = 8'b11000101;
DRAM[58552] = 8'b11001001;
DRAM[58553] = 8'b11010001;
DRAM[58554] = 8'b11011101;
DRAM[58555] = 8'b11101001;
DRAM[58556] = 8'b11110010;
DRAM[58557] = 8'b11110110;
DRAM[58558] = 8'b11110110;
DRAM[58559] = 8'b11110101;
DRAM[58560] = 8'b11111010;
DRAM[58561] = 8'b11110101;
DRAM[58562] = 8'b11011111;
DRAM[58563] = 8'b10111100;
DRAM[58564] = 8'b10100001;
DRAM[58565] = 8'b10010110;
DRAM[58566] = 8'b10010010;
DRAM[58567] = 8'b10001111;
DRAM[58568] = 8'b10001101;
DRAM[58569] = 8'b10001000;
DRAM[58570] = 8'b10000101;
DRAM[58571] = 8'b10001000;
DRAM[58572] = 8'b10001001;
DRAM[58573] = 8'b10000110;
DRAM[58574] = 8'b10000101;
DRAM[58575] = 8'b10000111;
DRAM[58576] = 8'b1111111;
DRAM[58577] = 8'b1111110;
DRAM[58578] = 8'b1111100;
DRAM[58579] = 8'b1111010;
DRAM[58580] = 8'b1111000;
DRAM[58581] = 8'b1110110;
DRAM[58582] = 8'b1110101;
DRAM[58583] = 8'b1110101;
DRAM[58584] = 8'b1110110;
DRAM[58585] = 8'b1110100;
DRAM[58586] = 8'b1110011;
DRAM[58587] = 8'b1110011;
DRAM[58588] = 8'b1110101;
DRAM[58589] = 8'b1110101;
DRAM[58590] = 8'b1110100;
DRAM[58591] = 8'b1110010;
DRAM[58592] = 8'b1101111;
DRAM[58593] = 8'b1101101;
DRAM[58594] = 8'b1101100;
DRAM[58595] = 8'b1101011;
DRAM[58596] = 8'b1101010;
DRAM[58597] = 8'b1101011;
DRAM[58598] = 8'b1101100;
DRAM[58599] = 8'b1101101;
DRAM[58600] = 8'b1101011;
DRAM[58601] = 8'b1101001;
DRAM[58602] = 8'b1100111;
DRAM[58603] = 8'b1100111;
DRAM[58604] = 8'b1101001;
DRAM[58605] = 8'b1101010;
DRAM[58606] = 8'b1101010;
DRAM[58607] = 8'b1101001;
DRAM[58608] = 8'b1101010;
DRAM[58609] = 8'b1101011;
DRAM[58610] = 8'b1101011;
DRAM[58611] = 8'b1101100;
DRAM[58612] = 8'b1101101;
DRAM[58613] = 8'b1101110;
DRAM[58614] = 8'b1101110;
DRAM[58615] = 8'b1101110;
DRAM[58616] = 8'b1101111;
DRAM[58617] = 8'b1101111;
DRAM[58618] = 8'b1101110;
DRAM[58619] = 8'b1101100;
DRAM[58620] = 8'b1101100;
DRAM[58621] = 8'b1101011;
DRAM[58622] = 8'b1101010;
DRAM[58623] = 8'b1101010;
DRAM[58624] = 8'b10001001;
DRAM[58625] = 8'b10001001;
DRAM[58626] = 8'b10001001;
DRAM[58627] = 8'b10001001;
DRAM[58628] = 8'b10001011;
DRAM[58629] = 8'b10001100;
DRAM[58630] = 8'b10001110;
DRAM[58631] = 8'b10001111;
DRAM[58632] = 8'b10010001;
DRAM[58633] = 8'b10010001;
DRAM[58634] = 8'b10010101;
DRAM[58635] = 8'b10011010;
DRAM[58636] = 8'b10100001;
DRAM[58637] = 8'b10110000;
DRAM[58638] = 8'b11001000;
DRAM[58639] = 8'b11011101;
DRAM[58640] = 8'b11110010;
DRAM[58641] = 8'b11110110;
DRAM[58642] = 8'b11111010;
DRAM[58643] = 8'b11111101;
DRAM[58644] = 8'b11111110;
DRAM[58645] = 8'b11111110;
DRAM[58646] = 8'b11111011;
DRAM[58647] = 8'b11111001;
DRAM[58648] = 8'b11111100;
DRAM[58649] = 8'b11110111;
DRAM[58650] = 8'b11110010;
DRAM[58651] = 8'b11101110;
DRAM[58652] = 8'b11101111;
DRAM[58653] = 8'b11110010;
DRAM[58654] = 8'b11110100;
DRAM[58655] = 8'b11110110;
DRAM[58656] = 8'b11110011;
DRAM[58657] = 8'b11110001;
DRAM[58658] = 8'b11101110;
DRAM[58659] = 8'b11101011;
DRAM[58660] = 8'b11100111;
DRAM[58661] = 8'b11100010;
DRAM[58662] = 8'b11011100;
DRAM[58663] = 8'b11011000;
DRAM[58664] = 8'b11010111;
DRAM[58665] = 8'b11010100;
DRAM[58666] = 8'b11010010;
DRAM[58667] = 8'b11010100;
DRAM[58668] = 8'b11010110;
DRAM[58669] = 8'b11010010;
DRAM[58670] = 8'b11001010;
DRAM[58671] = 8'b11000010;
DRAM[58672] = 8'b11000100;
DRAM[58673] = 8'b10110110;
DRAM[58674] = 8'b10111000;
DRAM[58675] = 8'b11001010;
DRAM[58676] = 8'b11001110;
DRAM[58677] = 8'b11000001;
DRAM[58678] = 8'b10111110;
DRAM[58679] = 8'b11001000;
DRAM[58680] = 8'b11000111;
DRAM[58681] = 8'b11001001;
DRAM[58682] = 8'b11001011;
DRAM[58683] = 8'b11001001;
DRAM[58684] = 8'b10111110;
DRAM[58685] = 8'b10110011;
DRAM[58686] = 8'b10110001;
DRAM[58687] = 8'b10110111;
DRAM[58688] = 8'b10110001;
DRAM[58689] = 8'b10110001;
DRAM[58690] = 8'b10101111;
DRAM[58691] = 8'b10101011;
DRAM[58692] = 8'b10100100;
DRAM[58693] = 8'b10011100;
DRAM[58694] = 8'b10010101;
DRAM[58695] = 8'b10010001;
DRAM[58696] = 8'b10010000;
DRAM[58697] = 8'b10001110;
DRAM[58698] = 8'b10001100;
DRAM[58699] = 8'b10001001;
DRAM[58700] = 8'b10000010;
DRAM[58701] = 8'b1111101;
DRAM[58702] = 8'b10000000;
DRAM[58703] = 8'b10001000;
DRAM[58704] = 8'b10000100;
DRAM[58705] = 8'b1110010;
DRAM[58706] = 8'b10000111;
DRAM[58707] = 8'b10010000;
DRAM[58708] = 8'b10000100;
DRAM[58709] = 8'b1111100;
DRAM[58710] = 8'b10001001;
DRAM[58711] = 8'b1111101;
DRAM[58712] = 8'b1110100;
DRAM[58713] = 8'b1110110;
DRAM[58714] = 8'b1111111;
DRAM[58715] = 8'b10000110;
DRAM[58716] = 8'b10000011;
DRAM[58717] = 8'b1111111;
DRAM[58718] = 8'b10001000;
DRAM[58719] = 8'b10010101;
DRAM[58720] = 8'b10000000;
DRAM[58721] = 8'b10000100;
DRAM[58722] = 8'b10000101;
DRAM[58723] = 8'b1111110;
DRAM[58724] = 8'b1111010;
DRAM[58725] = 8'b1111010;
DRAM[58726] = 8'b1111100;
DRAM[58727] = 8'b1111011;
DRAM[58728] = 8'b10000011;
DRAM[58729] = 8'b1110110;
DRAM[58730] = 8'b1110011;
DRAM[58731] = 8'b1110111;
DRAM[58732] = 8'b1110110;
DRAM[58733] = 8'b1111001;
DRAM[58734] = 8'b1111011;
DRAM[58735] = 8'b1110111;
DRAM[58736] = 8'b1101101;
DRAM[58737] = 8'b1100101;
DRAM[58738] = 8'b1101001;
DRAM[58739] = 8'b1101110;
DRAM[58740] = 8'b1101001;
DRAM[58741] = 8'b1101010;
DRAM[58742] = 8'b1101111;
DRAM[58743] = 8'b1101101;
DRAM[58744] = 8'b1110000;
DRAM[58745] = 8'b1110010;
DRAM[58746] = 8'b1110100;
DRAM[58747] = 8'b1110010;
DRAM[58748] = 8'b1101110;
DRAM[58749] = 8'b1101101;
DRAM[58750] = 8'b1101110;
DRAM[58751] = 8'b1110000;
DRAM[58752] = 8'b1101001;
DRAM[58753] = 8'b1110001;
DRAM[58754] = 8'b1110011;
DRAM[58755] = 8'b1101010;
DRAM[58756] = 8'b1100010;
DRAM[58757] = 8'b1100101;
DRAM[58758] = 8'b1101110;
DRAM[58759] = 8'b1110100;
DRAM[58760] = 8'b1101110;
DRAM[58761] = 8'b1101101;
DRAM[58762] = 8'b1101011;
DRAM[58763] = 8'b1101000;
DRAM[58764] = 8'b1101011;
DRAM[58765] = 8'b1101111;
DRAM[58766] = 8'b1101111;
DRAM[58767] = 8'b1101011;
DRAM[58768] = 8'b1100111;
DRAM[58769] = 8'b1101100;
DRAM[58770] = 8'b1101111;
DRAM[58771] = 8'b1101101;
DRAM[58772] = 8'b1101110;
DRAM[58773] = 8'b1110101;
DRAM[58774] = 8'b1111100;
DRAM[58775] = 8'b1111111;
DRAM[58776] = 8'b10000001;
DRAM[58777] = 8'b1110101;
DRAM[58778] = 8'b1110100;
DRAM[58779] = 8'b1111111;
DRAM[58780] = 8'b10000011;
DRAM[58781] = 8'b1111011;
DRAM[58782] = 8'b1110110;
DRAM[58783] = 8'b1111001;
DRAM[58784] = 8'b1111100;
DRAM[58785] = 8'b10000001;
DRAM[58786] = 8'b10000000;
DRAM[58787] = 8'b1111001;
DRAM[58788] = 8'b1110101;
DRAM[58789] = 8'b1111010;
DRAM[58790] = 8'b10000001;
DRAM[58791] = 8'b10000110;
DRAM[58792] = 8'b10001011;
DRAM[58793] = 8'b10010010;
DRAM[58794] = 8'b10010111;
DRAM[58795] = 8'b10011000;
DRAM[58796] = 8'b10011000;
DRAM[58797] = 8'b10011011;
DRAM[58798] = 8'b10011100;
DRAM[58799] = 8'b10011010;
DRAM[58800] = 8'b10100011;
DRAM[58801] = 8'b10100110;
DRAM[58802] = 8'b10101010;
DRAM[58803] = 8'b10101110;
DRAM[58804] = 8'b10110010;
DRAM[58805] = 8'b10111000;
DRAM[58806] = 8'b10111110;
DRAM[58807] = 8'b11000010;
DRAM[58808] = 8'b11000111;
DRAM[58809] = 8'b11001110;
DRAM[58810] = 8'b11011010;
DRAM[58811] = 8'b11100110;
DRAM[58812] = 8'b11101111;
DRAM[58813] = 8'b11110100;
DRAM[58814] = 8'b11110101;
DRAM[58815] = 8'b11110101;
DRAM[58816] = 8'b11111111;
DRAM[58817] = 8'b11111000;
DRAM[58818] = 8'b11100001;
DRAM[58819] = 8'b11000000;
DRAM[58820] = 8'b10100101;
DRAM[58821] = 8'b10011001;
DRAM[58822] = 8'b10010110;
DRAM[58823] = 8'b10010110;
DRAM[58824] = 8'b10010000;
DRAM[58825] = 8'b10001011;
DRAM[58826] = 8'b10001000;
DRAM[58827] = 8'b10001010;
DRAM[58828] = 8'b10001010;
DRAM[58829] = 8'b10000111;
DRAM[58830] = 8'b10000110;
DRAM[58831] = 8'b10000111;
DRAM[58832] = 8'b10000000;
DRAM[58833] = 8'b1111111;
DRAM[58834] = 8'b1111101;
DRAM[58835] = 8'b1111010;
DRAM[58836] = 8'b1111000;
DRAM[58837] = 8'b1110111;
DRAM[58838] = 8'b1110110;
DRAM[58839] = 8'b1110110;
DRAM[58840] = 8'b1110111;
DRAM[58841] = 8'b1110110;
DRAM[58842] = 8'b1110100;
DRAM[58843] = 8'b1110100;
DRAM[58844] = 8'b1110100;
DRAM[58845] = 8'b1110100;
DRAM[58846] = 8'b1110010;
DRAM[58847] = 8'b1110001;
DRAM[58848] = 8'b1101110;
DRAM[58849] = 8'b1101100;
DRAM[58850] = 8'b1101011;
DRAM[58851] = 8'b1101001;
DRAM[58852] = 8'b1101001;
DRAM[58853] = 8'b1101010;
DRAM[58854] = 8'b1101011;
DRAM[58855] = 8'b1101011;
DRAM[58856] = 8'b1101010;
DRAM[58857] = 8'b1101000;
DRAM[58858] = 8'b1100111;
DRAM[58859] = 8'b1100111;
DRAM[58860] = 8'b1101001;
DRAM[58861] = 8'b1101011;
DRAM[58862] = 8'b1101010;
DRAM[58863] = 8'b1101001;
DRAM[58864] = 8'b1101011;
DRAM[58865] = 8'b1101011;
DRAM[58866] = 8'b1101100;
DRAM[58867] = 8'b1101101;
DRAM[58868] = 8'b1101110;
DRAM[58869] = 8'b1101110;
DRAM[58870] = 8'b1101111;
DRAM[58871] = 8'b1101111;
DRAM[58872] = 8'b1110000;
DRAM[58873] = 8'b1101111;
DRAM[58874] = 8'b1101101;
DRAM[58875] = 8'b1101100;
DRAM[58876] = 8'b1101011;
DRAM[58877] = 8'b1101010;
DRAM[58878] = 8'b1101010;
DRAM[58879] = 8'b1101010;
DRAM[58880] = 8'b10001100;
DRAM[58881] = 8'b10001011;
DRAM[58882] = 8'b10001010;
DRAM[58883] = 8'b10001001;
DRAM[58884] = 8'b10001010;
DRAM[58885] = 8'b10001011;
DRAM[58886] = 8'b10001110;
DRAM[58887] = 8'b10001111;
DRAM[58888] = 8'b10010000;
DRAM[58889] = 8'b10001110;
DRAM[58890] = 8'b10010010;
DRAM[58891] = 8'b10011100;
DRAM[58892] = 8'b10101011;
DRAM[58893] = 8'b11000000;
DRAM[58894] = 8'b11011100;
DRAM[58895] = 8'b11110001;
DRAM[58896] = 8'b11111010;
DRAM[58897] = 8'b11111001;
DRAM[58898] = 8'b11111010;
DRAM[58899] = 8'b11111100;
DRAM[58900] = 8'b11111101;
DRAM[58901] = 8'b11111100;
DRAM[58902] = 8'b11111001;
DRAM[58903] = 8'b11110111;
DRAM[58904] = 8'b11111000;
DRAM[58905] = 8'b11110100;
DRAM[58906] = 8'b11110000;
DRAM[58907] = 8'b11101110;
DRAM[58908] = 8'b11101111;
DRAM[58909] = 8'b11110001;
DRAM[58910] = 8'b11110010;
DRAM[58911] = 8'b11110010;
DRAM[58912] = 8'b11101100;
DRAM[58913] = 8'b11101100;
DRAM[58914] = 8'b11101011;
DRAM[58915] = 8'b11100111;
DRAM[58916] = 8'b11100001;
DRAM[58917] = 8'b11011011;
DRAM[58918] = 8'b11010111;
DRAM[58919] = 8'b11010101;
DRAM[58920] = 8'b11010011;
DRAM[58921] = 8'b11010011;
DRAM[58922] = 8'b11010011;
DRAM[58923] = 8'b11010100;
DRAM[58924] = 8'b11010010;
DRAM[58925] = 8'b11001100;
DRAM[58926] = 8'b11000100;
DRAM[58927] = 8'b10111101;
DRAM[58928] = 8'b10111110;
DRAM[58929] = 8'b10101110;
DRAM[58930] = 8'b10101111;
DRAM[58931] = 8'b11000000;
DRAM[58932] = 8'b11000011;
DRAM[58933] = 8'b10110110;
DRAM[58934] = 8'b10111000;
DRAM[58935] = 8'b11001001;
DRAM[58936] = 8'b11000010;
DRAM[58937] = 8'b10110110;
DRAM[58938] = 8'b10101110;
DRAM[58939] = 8'b10110001;
DRAM[58940] = 8'b10111000;
DRAM[58941] = 8'b10110111;
DRAM[58942] = 8'b10110001;
DRAM[58943] = 8'b10101101;
DRAM[58944] = 8'b10100111;
DRAM[58945] = 8'b10101010;
DRAM[58946] = 8'b10101100;
DRAM[58947] = 8'b10101010;
DRAM[58948] = 8'b10100110;
DRAM[58949] = 8'b10100100;
DRAM[58950] = 8'b10100100;
DRAM[58951] = 8'b10100110;
DRAM[58952] = 8'b10011111;
DRAM[58953] = 8'b10010110;
DRAM[58954] = 8'b10001101;
DRAM[58955] = 8'b10000111;
DRAM[58956] = 8'b10000010;
DRAM[58957] = 8'b1111110;
DRAM[58958] = 8'b10000000;
DRAM[58959] = 8'b10000110;
DRAM[58960] = 8'b10000001;
DRAM[58961] = 8'b1110110;
DRAM[58962] = 8'b10000110;
DRAM[58963] = 8'b10011000;
DRAM[58964] = 8'b1111110;
DRAM[58965] = 8'b1111111;
DRAM[58966] = 8'b10000111;
DRAM[58967] = 8'b10000010;
DRAM[58968] = 8'b1111000;
DRAM[58969] = 8'b1110111;
DRAM[58970] = 8'b1111110;
DRAM[58971] = 8'b10000000;
DRAM[58972] = 8'b1111100;
DRAM[58973] = 8'b10000000;
DRAM[58974] = 8'b10001011;
DRAM[58975] = 8'b10010000;
DRAM[58976] = 8'b1111010;
DRAM[58977] = 8'b1111010;
DRAM[58978] = 8'b1111110;
DRAM[58979] = 8'b10000001;
DRAM[58980] = 8'b1111111;
DRAM[58981] = 8'b1111000;
DRAM[58982] = 8'b1110111;
DRAM[58983] = 8'b1111010;
DRAM[58984] = 8'b1111010;
DRAM[58985] = 8'b1111110;
DRAM[58986] = 8'b1111000;
DRAM[58987] = 8'b1110011;
DRAM[58988] = 8'b1111001;
DRAM[58989] = 8'b1111100;
DRAM[58990] = 8'b1111010;
DRAM[58991] = 8'b1111101;
DRAM[58992] = 8'b1110100;
DRAM[58993] = 8'b1101000;
DRAM[58994] = 8'b1101001;
DRAM[58995] = 8'b1110000;
DRAM[58996] = 8'b1101110;
DRAM[58997] = 8'b1101111;
DRAM[58998] = 8'b1110011;
DRAM[58999] = 8'b1110000;
DRAM[59000] = 8'b1110011;
DRAM[59001] = 8'b1110100;
DRAM[59002] = 8'b1110110;
DRAM[59003] = 8'b1110111;
DRAM[59004] = 8'b1110110;
DRAM[59005] = 8'b1110010;
DRAM[59006] = 8'b1110000;
DRAM[59007] = 8'b1110000;
DRAM[59008] = 8'b1101011;
DRAM[59009] = 8'b1101110;
DRAM[59010] = 8'b1110010;
DRAM[59011] = 8'b1110001;
DRAM[59012] = 8'b1101001;
DRAM[59013] = 8'b1100100;
DRAM[59014] = 8'b1101011;
DRAM[59015] = 8'b1110111;
DRAM[59016] = 8'b1110010;
DRAM[59017] = 8'b1110000;
DRAM[59018] = 8'b1101011;
DRAM[59019] = 8'b1101001;
DRAM[59020] = 8'b1101110;
DRAM[59021] = 8'b1110100;
DRAM[59022] = 8'b1110001;
DRAM[59023] = 8'b1101001;
DRAM[59024] = 8'b1110000;
DRAM[59025] = 8'b1101111;
DRAM[59026] = 8'b1110000;
DRAM[59027] = 8'b1110001;
DRAM[59028] = 8'b1110000;
DRAM[59029] = 8'b1101111;
DRAM[59030] = 8'b1110110;
DRAM[59031] = 8'b1111111;
DRAM[59032] = 8'b10000011;
DRAM[59033] = 8'b1110111;
DRAM[59034] = 8'b1110101;
DRAM[59035] = 8'b10000001;
DRAM[59036] = 8'b10000101;
DRAM[59037] = 8'b1111010;
DRAM[59038] = 8'b1110010;
DRAM[59039] = 8'b1110010;
DRAM[59040] = 8'b1110010;
DRAM[59041] = 8'b1111011;
DRAM[59042] = 8'b10000001;
DRAM[59043] = 8'b1111111;
DRAM[59044] = 8'b1111100;
DRAM[59045] = 8'b1111101;
DRAM[59046] = 8'b1111110;
DRAM[59047] = 8'b1111101;
DRAM[59048] = 8'b1111101;
DRAM[59049] = 8'b10001001;
DRAM[59050] = 8'b10010110;
DRAM[59051] = 8'b10011101;
DRAM[59052] = 8'b10011111;
DRAM[59053] = 8'b10011111;
DRAM[59054] = 8'b10011010;
DRAM[59055] = 8'b10010100;
DRAM[59056] = 8'b10011111;
DRAM[59057] = 8'b10100010;
DRAM[59058] = 8'b10101000;
DRAM[59059] = 8'b10101100;
DRAM[59060] = 8'b10110001;
DRAM[59061] = 8'b10110110;
DRAM[59062] = 8'b10111011;
DRAM[59063] = 8'b10111111;
DRAM[59064] = 8'b11001001;
DRAM[59065] = 8'b11001101;
DRAM[59066] = 8'b11010101;
DRAM[59067] = 8'b11011110;
DRAM[59068] = 8'b11100111;
DRAM[59069] = 8'b11101111;
DRAM[59070] = 8'b11110100;
DRAM[59071] = 8'b11110111;
DRAM[59072] = 8'b11111110;
DRAM[59073] = 8'b11111000;
DRAM[59074] = 8'b11100110;
DRAM[59075] = 8'b11001001;
DRAM[59076] = 8'b10101110;
DRAM[59077] = 8'b10011110;
DRAM[59078] = 8'b10010111;
DRAM[59079] = 8'b10010101;
DRAM[59080] = 8'b10010100;
DRAM[59081] = 8'b10001110;
DRAM[59082] = 8'b10001011;
DRAM[59083] = 8'b10001100;
DRAM[59084] = 8'b10001100;
DRAM[59085] = 8'b10001000;
DRAM[59086] = 8'b10000110;
DRAM[59087] = 8'b10000111;
DRAM[59088] = 8'b10000010;
DRAM[59089] = 8'b10000001;
DRAM[59090] = 8'b1111111;
DRAM[59091] = 8'b1111100;
DRAM[59092] = 8'b1111010;
DRAM[59093] = 8'b1111001;
DRAM[59094] = 8'b1111000;
DRAM[59095] = 8'b1111000;
DRAM[59096] = 8'b1111001;
DRAM[59097] = 8'b1110111;
DRAM[59098] = 8'b1110101;
DRAM[59099] = 8'b1110100;
DRAM[59100] = 8'b1110100;
DRAM[59101] = 8'b1110011;
DRAM[59102] = 8'b1110001;
DRAM[59103] = 8'b1101111;
DRAM[59104] = 8'b1101100;
DRAM[59105] = 8'b1101011;
DRAM[59106] = 8'b1101010;
DRAM[59107] = 8'b1101000;
DRAM[59108] = 8'b1101000;
DRAM[59109] = 8'b1101000;
DRAM[59110] = 8'b1101001;
DRAM[59111] = 8'b1101010;
DRAM[59112] = 8'b1101010;
DRAM[59113] = 8'b1101000;
DRAM[59114] = 8'b1100111;
DRAM[59115] = 8'b1100111;
DRAM[59116] = 8'b1101001;
DRAM[59117] = 8'b1101011;
DRAM[59118] = 8'b1101011;
DRAM[59119] = 8'b1101010;
DRAM[59120] = 8'b1101100;
DRAM[59121] = 8'b1101100;
DRAM[59122] = 8'b1101101;
DRAM[59123] = 8'b1101101;
DRAM[59124] = 8'b1101110;
DRAM[59125] = 8'b1101111;
DRAM[59126] = 8'b1110000;
DRAM[59127] = 8'b1110000;
DRAM[59128] = 8'b1110000;
DRAM[59129] = 8'b1101111;
DRAM[59130] = 8'b1101101;
DRAM[59131] = 8'b1101011;
DRAM[59132] = 8'b1101001;
DRAM[59133] = 8'b1101001;
DRAM[59134] = 8'b1101001;
DRAM[59135] = 8'b1101001;
DRAM[59136] = 8'b10001111;
DRAM[59137] = 8'b10001101;
DRAM[59138] = 8'b10001010;
DRAM[59139] = 8'b10001001;
DRAM[59140] = 8'b10001001;
DRAM[59141] = 8'b10001011;
DRAM[59142] = 8'b10001110;
DRAM[59143] = 8'b10010000;
DRAM[59144] = 8'b10010000;
DRAM[59145] = 8'b10001101;
DRAM[59146] = 8'b10010000;
DRAM[59147] = 8'b10011101;
DRAM[59148] = 8'b10101111;
DRAM[59149] = 8'b11001000;
DRAM[59150] = 8'b11100100;
DRAM[59151] = 8'b11111001;
DRAM[59152] = 8'b11111010;
DRAM[59153] = 8'b11110111;
DRAM[59154] = 8'b11110110;
DRAM[59155] = 8'b11111001;
DRAM[59156] = 8'b11111100;
DRAM[59157] = 8'b11111011;
DRAM[59158] = 8'b11111000;
DRAM[59159] = 8'b11110111;
DRAM[59160] = 8'b11110100;
DRAM[59161] = 8'b11110001;
DRAM[59162] = 8'b11101111;
DRAM[59163] = 8'b11101110;
DRAM[59164] = 8'b11101110;
DRAM[59165] = 8'b11101110;
DRAM[59166] = 8'b11101101;
DRAM[59167] = 8'b11101100;
DRAM[59168] = 8'b11100111;
DRAM[59169] = 8'b11101010;
DRAM[59170] = 8'b11101011;
DRAM[59171] = 8'b11101000;
DRAM[59172] = 8'b11100010;
DRAM[59173] = 8'b11011110;
DRAM[59174] = 8'b11011100;
DRAM[59175] = 8'b11011101;
DRAM[59176] = 8'b11010000;
DRAM[59177] = 8'b11010001;
DRAM[59178] = 8'b11010011;
DRAM[59179] = 8'b11010010;
DRAM[59180] = 8'b11001110;
DRAM[59181] = 8'b11000110;
DRAM[59182] = 8'b10111111;
DRAM[59183] = 8'b10111010;
DRAM[59184] = 8'b10110010;
DRAM[59185] = 8'b10110010;
DRAM[59186] = 8'b10110000;
DRAM[59187] = 8'b10101101;
DRAM[59188] = 8'b10101101;
DRAM[59189] = 8'b10110001;
DRAM[59190] = 8'b10110111;
DRAM[59191] = 8'b10111010;
DRAM[59192] = 8'b10111010;
DRAM[59193] = 8'b10110100;
DRAM[59194] = 8'b10101111;
DRAM[59195] = 8'b10101100;
DRAM[59196] = 8'b10100110;
DRAM[59197] = 8'b10100010;
DRAM[59198] = 8'b10100100;
DRAM[59199] = 8'b10101010;
DRAM[59200] = 8'b10100010;
DRAM[59201] = 8'b10100101;
DRAM[59202] = 8'b10100111;
DRAM[59203] = 8'b10100100;
DRAM[59204] = 8'b10011111;
DRAM[59205] = 8'b10011110;
DRAM[59206] = 8'b10100011;
DRAM[59207] = 8'b10101001;
DRAM[59208] = 8'b10011101;
DRAM[59209] = 8'b10010010;
DRAM[59210] = 8'b10001010;
DRAM[59211] = 8'b10001011;
DRAM[59212] = 8'b10001111;
DRAM[59213] = 8'b10001111;
DRAM[59214] = 8'b10001111;
DRAM[59215] = 8'b10010000;
DRAM[59216] = 8'b1111100;
DRAM[59217] = 8'b10010000;
DRAM[59218] = 8'b1111111;
DRAM[59219] = 8'b10000111;
DRAM[59220] = 8'b10000100;
DRAM[59221] = 8'b10000010;
DRAM[59222] = 8'b1110100;
DRAM[59223] = 8'b10010110;
DRAM[59224] = 8'b10000110;
DRAM[59225] = 8'b10000000;
DRAM[59226] = 8'b10000001;
DRAM[59227] = 8'b1111110;
DRAM[59228] = 8'b1111000;
DRAM[59229] = 8'b10000000;
DRAM[59230] = 8'b10001011;
DRAM[59231] = 8'b10001000;
DRAM[59232] = 8'b1111001;
DRAM[59233] = 8'b1110011;
DRAM[59234] = 8'b1110111;
DRAM[59235] = 8'b10000010;
DRAM[59236] = 8'b10000011;
DRAM[59237] = 8'b1111000;
DRAM[59238] = 8'b1110100;
DRAM[59239] = 8'b1111001;
DRAM[59240] = 8'b1110111;
DRAM[59241] = 8'b10000111;
DRAM[59242] = 8'b1111101;
DRAM[59243] = 8'b1110000;
DRAM[59244] = 8'b1111001;
DRAM[59245] = 8'b1111100;
DRAM[59246] = 8'b1110110;
DRAM[59247] = 8'b1111100;
DRAM[59248] = 8'b1111011;
DRAM[59249] = 8'b1101011;
DRAM[59250] = 8'b1101001;
DRAM[59251] = 8'b1110000;
DRAM[59252] = 8'b1110000;
DRAM[59253] = 8'b1110010;
DRAM[59254] = 8'b1110111;
DRAM[59255] = 8'b1110100;
DRAM[59256] = 8'b1110010;
DRAM[59257] = 8'b1110011;
DRAM[59258] = 8'b1110110;
DRAM[59259] = 8'b1111011;
DRAM[59260] = 8'b1111010;
DRAM[59261] = 8'b1110101;
DRAM[59262] = 8'b1110000;
DRAM[59263] = 8'b1101110;
DRAM[59264] = 8'b1101100;
DRAM[59265] = 8'b1101100;
DRAM[59266] = 8'b1110010;
DRAM[59267] = 8'b1110111;
DRAM[59268] = 8'b1110000;
DRAM[59269] = 8'b1100101;
DRAM[59270] = 8'b1101010;
DRAM[59271] = 8'b1111001;
DRAM[59272] = 8'b1110110;
DRAM[59273] = 8'b1110000;
DRAM[59274] = 8'b1100111;
DRAM[59275] = 8'b1100101;
DRAM[59276] = 8'b1101111;
DRAM[59277] = 8'b1111000;
DRAM[59278] = 8'b1110010;
DRAM[59279] = 8'b1100110;
DRAM[59280] = 8'b1111010;
DRAM[59281] = 8'b1110101;
DRAM[59282] = 8'b1110100;
DRAM[59283] = 8'b1110101;
DRAM[59284] = 8'b1110000;
DRAM[59285] = 8'b1101001;
DRAM[59286] = 8'b1101110;
DRAM[59287] = 8'b1111010;
DRAM[59288] = 8'b1110100;
DRAM[59289] = 8'b1111010;
DRAM[59290] = 8'b1111011;
DRAM[59291] = 8'b1111000;
DRAM[59292] = 8'b1111110;
DRAM[59293] = 8'b10000110;
DRAM[59294] = 8'b1111101;
DRAM[59295] = 8'b1101100;
DRAM[59296] = 8'b1101111;
DRAM[59297] = 8'b1111000;
DRAM[59298] = 8'b10000000;
DRAM[59299] = 8'b10000011;
DRAM[59300] = 8'b10000101;
DRAM[59301] = 8'b10001000;
DRAM[59302] = 8'b10000110;
DRAM[59303] = 8'b10000010;
DRAM[59304] = 8'b10000101;
DRAM[59305] = 8'b10001000;
DRAM[59306] = 8'b10001001;
DRAM[59307] = 8'b10001000;
DRAM[59308] = 8'b10001100;
DRAM[59309] = 8'b10010111;
DRAM[59310] = 8'b10100000;
DRAM[59311] = 8'b10100100;
DRAM[59312] = 8'b10011010;
DRAM[59313] = 8'b10011111;
DRAM[59314] = 8'b10100110;
DRAM[59315] = 8'b10101101;
DRAM[59316] = 8'b10110011;
DRAM[59317] = 8'b10111001;
DRAM[59318] = 8'b10111111;
DRAM[59319] = 8'b11000011;
DRAM[59320] = 8'b11010000;
DRAM[59321] = 8'b11010010;
DRAM[59322] = 8'b11010110;
DRAM[59323] = 8'b11011100;
DRAM[59324] = 8'b11100110;
DRAM[59325] = 8'b11110000;
DRAM[59326] = 8'b11111001;
DRAM[59327] = 8'b11111110;
DRAM[59328] = 8'b11111000;
DRAM[59329] = 8'b11110101;
DRAM[59330] = 8'b11101001;
DRAM[59331] = 8'b11010000;
DRAM[59332] = 8'b10110101;
DRAM[59333] = 8'b10100001;
DRAM[59334] = 8'b10010101;
DRAM[59335] = 8'b10010000;
DRAM[59336] = 8'b10010110;
DRAM[59337] = 8'b10010000;
DRAM[59338] = 8'b10001101;
DRAM[59339] = 8'b10001101;
DRAM[59340] = 8'b10001100;
DRAM[59341] = 8'b10001000;
DRAM[59342] = 8'b10000110;
DRAM[59343] = 8'b10000111;
DRAM[59344] = 8'b10000100;
DRAM[59345] = 8'b10000011;
DRAM[59346] = 8'b10000001;
DRAM[59347] = 8'b1111110;
DRAM[59348] = 8'b1111100;
DRAM[59349] = 8'b1111011;
DRAM[59350] = 8'b1111010;
DRAM[59351] = 8'b1111010;
DRAM[59352] = 8'b1111010;
DRAM[59353] = 8'b1111000;
DRAM[59354] = 8'b1110110;
DRAM[59355] = 8'b1110100;
DRAM[59356] = 8'b1110100;
DRAM[59357] = 8'b1110010;
DRAM[59358] = 8'b1110000;
DRAM[59359] = 8'b1101110;
DRAM[59360] = 8'b1101011;
DRAM[59361] = 8'b1101010;
DRAM[59362] = 8'b1101001;
DRAM[59363] = 8'b1100111;
DRAM[59364] = 8'b1100111;
DRAM[59365] = 8'b1101000;
DRAM[59366] = 8'b1101001;
DRAM[59367] = 8'b1101001;
DRAM[59368] = 8'b1101010;
DRAM[59369] = 8'b1101000;
DRAM[59370] = 8'b1100110;
DRAM[59371] = 8'b1100111;
DRAM[59372] = 8'b1101001;
DRAM[59373] = 8'b1101011;
DRAM[59374] = 8'b1101011;
DRAM[59375] = 8'b1101010;
DRAM[59376] = 8'b1101100;
DRAM[59377] = 8'b1101100;
DRAM[59378] = 8'b1101101;
DRAM[59379] = 8'b1101110;
DRAM[59380] = 8'b1101111;
DRAM[59381] = 8'b1101111;
DRAM[59382] = 8'b1110000;
DRAM[59383] = 8'b1110000;
DRAM[59384] = 8'b1110000;
DRAM[59385] = 8'b1101111;
DRAM[59386] = 8'b1101100;
DRAM[59387] = 8'b1101010;
DRAM[59388] = 8'b1101001;
DRAM[59389] = 8'b1101000;
DRAM[59390] = 8'b1101001;
DRAM[59391] = 8'b1101001;
DRAM[59392] = 8'b10001111;
DRAM[59393] = 8'b10001110;
DRAM[59394] = 8'b10001101;
DRAM[59395] = 8'b10001100;
DRAM[59396] = 8'b10001100;
DRAM[59397] = 8'b10001011;
DRAM[59398] = 8'b10001100;
DRAM[59399] = 8'b10001100;
DRAM[59400] = 8'b10001010;
DRAM[59401] = 8'b10010100;
DRAM[59402] = 8'b10011010;
DRAM[59403] = 8'b10011111;
DRAM[59404] = 8'b10110011;
DRAM[59405] = 8'b11010101;
DRAM[59406] = 8'b11101111;
DRAM[59407] = 8'b11111000;
DRAM[59408] = 8'b11110110;
DRAM[59409] = 8'b11111001;
DRAM[59410] = 8'b11111100;
DRAM[59411] = 8'b11111110;
DRAM[59412] = 8'b11111101;
DRAM[59413] = 8'b11111011;
DRAM[59414] = 8'b11111001;
DRAM[59415] = 8'b11111000;
DRAM[59416] = 8'b11110000;
DRAM[59417] = 8'b11101111;
DRAM[59418] = 8'b11101111;
DRAM[59419] = 8'b11110001;
DRAM[59420] = 8'b11110010;
DRAM[59421] = 8'b11110010;
DRAM[59422] = 8'b11110000;
DRAM[59423] = 8'b11101110;
DRAM[59424] = 8'b11101100;
DRAM[59425] = 8'b11100111;
DRAM[59426] = 8'b11100000;
DRAM[59427] = 8'b11011100;
DRAM[59428] = 8'b11011010;
DRAM[59429] = 8'b11011001;
DRAM[59430] = 8'b11011001;
DRAM[59431] = 8'b11011000;
DRAM[59432] = 8'b11011011;
DRAM[59433] = 8'b11011010;
DRAM[59434] = 8'b11010111;
DRAM[59435] = 8'b11010010;
DRAM[59436] = 8'b11001100;
DRAM[59437] = 8'b11000101;
DRAM[59438] = 8'b10111111;
DRAM[59439] = 8'b10111100;
DRAM[59440] = 8'b10110110;
DRAM[59441] = 8'b10101101;
DRAM[59442] = 8'b10100100;
DRAM[59443] = 8'b10100011;
DRAM[59444] = 8'b10101000;
DRAM[59445] = 8'b10101100;
DRAM[59446] = 8'b10101100;
DRAM[59447] = 8'b10101001;
DRAM[59448] = 8'b10100000;
DRAM[59449] = 8'b10100101;
DRAM[59450] = 8'b10100110;
DRAM[59451] = 8'b10100011;
DRAM[59452] = 8'b10100100;
DRAM[59453] = 8'b10101000;
DRAM[59454] = 8'b10101000;
DRAM[59455] = 8'b10100100;
DRAM[59456] = 8'b10100001;
DRAM[59457] = 8'b10101000;
DRAM[59458] = 8'b10100011;
DRAM[59459] = 8'b10011000;
DRAM[59460] = 8'b10011110;
DRAM[59461] = 8'b10101111;
DRAM[59462] = 8'b10110100;
DRAM[59463] = 8'b10101011;
DRAM[59464] = 8'b10010111;
DRAM[59465] = 8'b10010100;
DRAM[59466] = 8'b10011010;
DRAM[59467] = 8'b10010001;
DRAM[59468] = 8'b10000000;
DRAM[59469] = 8'b10001011;
DRAM[59470] = 8'b10011000;
DRAM[59471] = 8'b10001100;
DRAM[59472] = 8'b1111101;
DRAM[59473] = 8'b10000000;
DRAM[59474] = 8'b10001010;
DRAM[59475] = 8'b10000110;
DRAM[59476] = 8'b1111101;
DRAM[59477] = 8'b10001110;
DRAM[59478] = 8'b10010010;
DRAM[59479] = 8'b1111000;
DRAM[59480] = 8'b1111000;
DRAM[59481] = 8'b10001001;
DRAM[59482] = 8'b1101111;
DRAM[59483] = 8'b1101100;
DRAM[59484] = 8'b1101110;
DRAM[59485] = 8'b1101011;
DRAM[59486] = 8'b10000101;
DRAM[59487] = 8'b10001001;
DRAM[59488] = 8'b1110001;
DRAM[59489] = 8'b1110000;
DRAM[59490] = 8'b1111101;
DRAM[59491] = 8'b1111001;
DRAM[59492] = 8'b1111101;
DRAM[59493] = 8'b10000011;
DRAM[59494] = 8'b1110000;
DRAM[59495] = 8'b1101001;
DRAM[59496] = 8'b1110110;
DRAM[59497] = 8'b1111100;
DRAM[59498] = 8'b1111101;
DRAM[59499] = 8'b1110111;
DRAM[59500] = 8'b1110101;
DRAM[59501] = 8'b1111001;
DRAM[59502] = 8'b1111100;
DRAM[59503] = 8'b1111011;
DRAM[59504] = 8'b1111001;
DRAM[59505] = 8'b1110101;
DRAM[59506] = 8'b1110000;
DRAM[59507] = 8'b1101101;
DRAM[59508] = 8'b1101110;
DRAM[59509] = 8'b1110011;
DRAM[59510] = 8'b1111000;
DRAM[59511] = 8'b1111011;
DRAM[59512] = 8'b1100111;
DRAM[59513] = 8'b1111111;
DRAM[59514] = 8'b1110110;
DRAM[59515] = 8'b1110011;
DRAM[59516] = 8'b1111010;
DRAM[59517] = 8'b1111010;
DRAM[59518] = 8'b1110111;
DRAM[59519] = 8'b1100110;
DRAM[59520] = 8'b1101011;
DRAM[59521] = 8'b1101001;
DRAM[59522] = 8'b1110010;
DRAM[59523] = 8'b1100111;
DRAM[59524] = 8'b1100101;
DRAM[59525] = 8'b1101111;
DRAM[59526] = 8'b1101011;
DRAM[59527] = 8'b1110010;
DRAM[59528] = 8'b1110010;
DRAM[59529] = 8'b1101100;
DRAM[59530] = 8'b1101000;
DRAM[59531] = 8'b1101100;
DRAM[59532] = 8'b1101111;
DRAM[59533] = 8'b1101111;
DRAM[59534] = 8'b1101100;
DRAM[59535] = 8'b1101010;
DRAM[59536] = 8'b1101000;
DRAM[59537] = 8'b1111000;
DRAM[59538] = 8'b1101100;
DRAM[59539] = 8'b1100111;
DRAM[59540] = 8'b1111010;
DRAM[59541] = 8'b1110110;
DRAM[59542] = 8'b1101011;
DRAM[59543] = 8'b1111011;
DRAM[59544] = 8'b1110101;
DRAM[59545] = 8'b1111001;
DRAM[59546] = 8'b1110111;
DRAM[59547] = 8'b1110010;
DRAM[59548] = 8'b1111000;
DRAM[59549] = 8'b10000000;
DRAM[59550] = 8'b1111011;
DRAM[59551] = 8'b1101110;
DRAM[59552] = 8'b1110110;
DRAM[59553] = 8'b1110010;
DRAM[59554] = 8'b1111110;
DRAM[59555] = 8'b1111100;
DRAM[59556] = 8'b1111111;
DRAM[59557] = 8'b10001000;
DRAM[59558] = 8'b10000011;
DRAM[59559] = 8'b10001011;
DRAM[59560] = 8'b10000010;
DRAM[59561] = 8'b10000000;
DRAM[59562] = 8'b10000000;
DRAM[59563] = 8'b10000100;
DRAM[59564] = 8'b10001100;
DRAM[59565] = 8'b10010100;
DRAM[59566] = 8'b10011010;
DRAM[59567] = 8'b10011101;
DRAM[59568] = 8'b10011111;
DRAM[59569] = 8'b10100000;
DRAM[59570] = 8'b10100111;
DRAM[59571] = 8'b10101111;
DRAM[59572] = 8'b10110100;
DRAM[59573] = 8'b10110110;
DRAM[59574] = 8'b10111011;
DRAM[59575] = 8'b11000001;
DRAM[59576] = 8'b11001101;
DRAM[59577] = 8'b11010000;
DRAM[59578] = 8'b11010101;
DRAM[59579] = 8'b11011111;
DRAM[59580] = 8'b11101001;
DRAM[59581] = 8'b11110001;
DRAM[59582] = 8'b11110110;
DRAM[59583] = 8'b11110111;
DRAM[59584] = 8'b11110010;
DRAM[59585] = 8'b11110100;
DRAM[59586] = 8'b11100111;
DRAM[59587] = 8'b11001001;
DRAM[59588] = 8'b10110001;
DRAM[59589] = 8'b10100110;
DRAM[59590] = 8'b10011110;
DRAM[59591] = 8'b10010101;
DRAM[59592] = 8'b10001110;
DRAM[59593] = 8'b10001110;
DRAM[59594] = 8'b10001110;
DRAM[59595] = 8'b10001101;
DRAM[59596] = 8'b10001100;
DRAM[59597] = 8'b10001011;
DRAM[59598] = 8'b10001001;
DRAM[59599] = 8'b10001001;
DRAM[59600] = 8'b10000001;
DRAM[59601] = 8'b10000001;
DRAM[59602] = 8'b1111111;
DRAM[59603] = 8'b1111101;
DRAM[59604] = 8'b1111011;
DRAM[59605] = 8'b1111001;
DRAM[59606] = 8'b1111000;
DRAM[59607] = 8'b1110111;
DRAM[59608] = 8'b1110110;
DRAM[59609] = 8'b1110110;
DRAM[59610] = 8'b1110101;
DRAM[59611] = 8'b1110011;
DRAM[59612] = 8'b1110001;
DRAM[59613] = 8'b1101111;
DRAM[59614] = 8'b1101110;
DRAM[59615] = 8'b1101101;
DRAM[59616] = 8'b1101100;
DRAM[59617] = 8'b1101011;
DRAM[59618] = 8'b1101010;
DRAM[59619] = 8'b1101001;
DRAM[59620] = 8'b1101001;
DRAM[59621] = 8'b1101001;
DRAM[59622] = 8'b1101001;
DRAM[59623] = 8'b1101010;
DRAM[59624] = 8'b1101000;
DRAM[59625] = 8'b1100111;
DRAM[59626] = 8'b1100111;
DRAM[59627] = 8'b1100111;
DRAM[59628] = 8'b1100111;
DRAM[59629] = 8'b1101000;
DRAM[59630] = 8'b1101001;
DRAM[59631] = 8'b1101010;
DRAM[59632] = 8'b1101101;
DRAM[59633] = 8'b1101100;
DRAM[59634] = 8'b1101011;
DRAM[59635] = 8'b1101101;
DRAM[59636] = 8'b1101111;
DRAM[59637] = 8'b1110001;
DRAM[59638] = 8'b1110000;
DRAM[59639] = 8'b1101111;
DRAM[59640] = 8'b1101100;
DRAM[59641] = 8'b1101100;
DRAM[59642] = 8'b1101100;
DRAM[59643] = 8'b1101011;
DRAM[59644] = 8'b1101010;
DRAM[59645] = 8'b1101001;
DRAM[59646] = 8'b1100111;
DRAM[59647] = 8'b1100110;
DRAM[59648] = 8'b10010011;
DRAM[59649] = 8'b10010010;
DRAM[59650] = 8'b10010000;
DRAM[59651] = 8'b10001111;
DRAM[59652] = 8'b10001110;
DRAM[59653] = 8'b10001110;
DRAM[59654] = 8'b10001111;
DRAM[59655] = 8'b10001111;
DRAM[59656] = 8'b10000111;
DRAM[59657] = 8'b10001111;
DRAM[59658] = 8'b10010110;
DRAM[59659] = 8'b10011110;
DRAM[59660] = 8'b10110111;
DRAM[59661] = 8'b11011010;
DRAM[59662] = 8'b11110010;
DRAM[59663] = 8'b11111001;
DRAM[59664] = 8'b11111001;
DRAM[59665] = 8'b11111011;
DRAM[59666] = 8'b11111101;
DRAM[59667] = 8'b11111110;
DRAM[59668] = 8'b11111100;
DRAM[59669] = 8'b11111001;
DRAM[59670] = 8'b11110110;
DRAM[59671] = 8'b11110101;
DRAM[59672] = 8'b11110100;
DRAM[59673] = 8'b11110001;
DRAM[59674] = 8'b11101111;
DRAM[59675] = 8'b11101101;
DRAM[59676] = 8'b11101110;
DRAM[59677] = 8'b11101110;
DRAM[59678] = 8'b11101100;
DRAM[59679] = 8'b11101011;
DRAM[59680] = 8'b11100010;
DRAM[59681] = 8'b11100000;
DRAM[59682] = 8'b11011101;
DRAM[59683] = 8'b11011100;
DRAM[59684] = 8'b11011010;
DRAM[59685] = 8'b11010111;
DRAM[59686] = 8'b11010010;
DRAM[59687] = 8'b11001110;
DRAM[59688] = 8'b11010010;
DRAM[59689] = 8'b11010010;
DRAM[59690] = 8'b11010000;
DRAM[59691] = 8'b11001100;
DRAM[59692] = 8'b11001000;
DRAM[59693] = 8'b11000011;
DRAM[59694] = 8'b10111111;
DRAM[59695] = 8'b10111100;
DRAM[59696] = 8'b10111011;
DRAM[59697] = 8'b10110010;
DRAM[59698] = 8'b10100111;
DRAM[59699] = 8'b10100010;
DRAM[59700] = 8'b10100001;
DRAM[59701] = 8'b10011110;
DRAM[59702] = 8'b10011000;
DRAM[59703] = 8'b10010010;
DRAM[59704] = 8'b10010011;
DRAM[59705] = 8'b10100001;
DRAM[59706] = 8'b10101001;
DRAM[59707] = 8'b10100000;
DRAM[59708] = 8'b10010100;
DRAM[59709] = 8'b10010010;
DRAM[59710] = 8'b10011001;
DRAM[59711] = 8'b10011111;
DRAM[59712] = 8'b10010100;
DRAM[59713] = 8'b10011001;
DRAM[59714] = 8'b10011010;
DRAM[59715] = 8'b10011011;
DRAM[59716] = 8'b10100100;
DRAM[59717] = 8'b10101101;
DRAM[59718] = 8'b10101000;
DRAM[59719] = 8'b10011011;
DRAM[59720] = 8'b10011100;
DRAM[59721] = 8'b10011000;
DRAM[59722] = 8'b10010101;
DRAM[59723] = 8'b10010000;
DRAM[59724] = 8'b10010000;
DRAM[59725] = 8'b10011001;
DRAM[59726] = 8'b10010111;
DRAM[59727] = 8'b10000110;
DRAM[59728] = 8'b1111101;
DRAM[59729] = 8'b1111100;
DRAM[59730] = 8'b10000001;
DRAM[59731] = 8'b10000011;
DRAM[59732] = 8'b10000000;
DRAM[59733] = 8'b10000011;
DRAM[59734] = 8'b10000101;
DRAM[59735] = 8'b1111101;
DRAM[59736] = 8'b1111100;
DRAM[59737] = 8'b10000100;
DRAM[59738] = 8'b1110011;
DRAM[59739] = 8'b1101101;
DRAM[59740] = 8'b1110010;
DRAM[59741] = 8'b1110010;
DRAM[59742] = 8'b1111001;
DRAM[59743] = 8'b1111011;
DRAM[59744] = 8'b10000010;
DRAM[59745] = 8'b1110110;
DRAM[59746] = 8'b1111010;
DRAM[59747] = 8'b1110110;
DRAM[59748] = 8'b1111001;
DRAM[59749] = 8'b1111110;
DRAM[59750] = 8'b1110011;
DRAM[59751] = 8'b1110111;
DRAM[59752] = 8'b1100111;
DRAM[59753] = 8'b1110110;
DRAM[59754] = 8'b10000000;
DRAM[59755] = 8'b1111010;
DRAM[59756] = 8'b1101111;
DRAM[59757] = 8'b1101111;
DRAM[59758] = 8'b1110111;
DRAM[59759] = 8'b1111110;
DRAM[59760] = 8'b1100011;
DRAM[59761] = 8'b1110010;
DRAM[59762] = 8'b10000000;
DRAM[59763] = 8'b10000000;
DRAM[59764] = 8'b1110101;
DRAM[59765] = 8'b1101110;
DRAM[59766] = 8'b1110100;
DRAM[59767] = 8'b1111101;
DRAM[59768] = 8'b1110010;
DRAM[59769] = 8'b10000011;
DRAM[59770] = 8'b1110110;
DRAM[59771] = 8'b1110100;
DRAM[59772] = 8'b1111010;
DRAM[59773] = 8'b1110101;
DRAM[59774] = 8'b1110100;
DRAM[59775] = 8'b1101000;
DRAM[59776] = 8'b1101111;
DRAM[59777] = 8'b1101010;
DRAM[59778] = 8'b1110010;
DRAM[59779] = 8'b1101011;
DRAM[59780] = 8'b1101010;
DRAM[59781] = 8'b1110000;
DRAM[59782] = 8'b1101100;
DRAM[59783] = 8'b1110110;
DRAM[59784] = 8'b1111000;
DRAM[59785] = 8'b1110011;
DRAM[59786] = 8'b1101101;
DRAM[59787] = 8'b1101011;
DRAM[59788] = 8'b1101111;
DRAM[59789] = 8'b1110011;
DRAM[59790] = 8'b1110011;
DRAM[59791] = 8'b1110000;
DRAM[59792] = 8'b1100010;
DRAM[59793] = 8'b1110001;
DRAM[59794] = 8'b1101111;
DRAM[59795] = 8'b1101110;
DRAM[59796] = 8'b1111000;
DRAM[59797] = 8'b1110101;
DRAM[59798] = 8'b1110000;
DRAM[59799] = 8'b1111101;
DRAM[59800] = 8'b1111100;
DRAM[59801] = 8'b1110011;
DRAM[59802] = 8'b1100111;
DRAM[59803] = 8'b1101001;
DRAM[59804] = 8'b1111100;
DRAM[59805] = 8'b10001011;
DRAM[59806] = 8'b1111110;
DRAM[59807] = 8'b1100111;
DRAM[59808] = 8'b1110001;
DRAM[59809] = 8'b1101100;
DRAM[59810] = 8'b1110110;
DRAM[59811] = 8'b1110001;
DRAM[59812] = 8'b1110001;
DRAM[59813] = 8'b1111000;
DRAM[59814] = 8'b1110010;
DRAM[59815] = 8'b1111001;
DRAM[59816] = 8'b10000110;
DRAM[59817] = 8'b10000101;
DRAM[59818] = 8'b10000100;
DRAM[59819] = 8'b10000001;
DRAM[59820] = 8'b1111111;
DRAM[59821] = 8'b10000010;
DRAM[59822] = 8'b10001000;
DRAM[59823] = 8'b10001101;
DRAM[59824] = 8'b10011111;
DRAM[59825] = 8'b10100000;
DRAM[59826] = 8'b10100101;
DRAM[59827] = 8'b10101101;
DRAM[59828] = 8'b10110001;
DRAM[59829] = 8'b10110011;
DRAM[59830] = 8'b10111001;
DRAM[59831] = 8'b10111111;
DRAM[59832] = 8'b11001010;
DRAM[59833] = 8'b11001110;
DRAM[59834] = 8'b11010100;
DRAM[59835] = 8'b11011101;
DRAM[59836] = 8'b11100101;
DRAM[59837] = 8'b11101101;
DRAM[59838] = 8'b11110100;
DRAM[59839] = 8'b11110111;
DRAM[59840] = 8'b11111000;
DRAM[59841] = 8'b11110110;
DRAM[59842] = 8'b11100010;
DRAM[59843] = 8'b10111111;
DRAM[59844] = 8'b10100100;
DRAM[59845] = 8'b10011011;
DRAM[59846] = 8'b10011001;
DRAM[59847] = 8'b10010110;
DRAM[59848] = 8'b10010001;
DRAM[59849] = 8'b10010000;
DRAM[59850] = 8'b10001111;
DRAM[59851] = 8'b10001110;
DRAM[59852] = 8'b10001100;
DRAM[59853] = 8'b10001001;
DRAM[59854] = 8'b10000111;
DRAM[59855] = 8'b10000110;
DRAM[59856] = 8'b10000000;
DRAM[59857] = 8'b1111111;
DRAM[59858] = 8'b1111101;
DRAM[59859] = 8'b1111010;
DRAM[59860] = 8'b1111000;
DRAM[59861] = 8'b1110111;
DRAM[59862] = 8'b1110110;
DRAM[59863] = 8'b1110110;
DRAM[59864] = 8'b1110111;
DRAM[59865] = 8'b1110110;
DRAM[59866] = 8'b1110101;
DRAM[59867] = 8'b1110011;
DRAM[59868] = 8'b1110001;
DRAM[59869] = 8'b1110000;
DRAM[59870] = 8'b1101111;
DRAM[59871] = 8'b1101110;
DRAM[59872] = 8'b1101100;
DRAM[59873] = 8'b1101011;
DRAM[59874] = 8'b1101010;
DRAM[59875] = 8'b1101001;
DRAM[59876] = 8'b1101001;
DRAM[59877] = 8'b1101001;
DRAM[59878] = 8'b1101001;
DRAM[59879] = 8'b1101010;
DRAM[59880] = 8'b1101000;
DRAM[59881] = 8'b1100111;
DRAM[59882] = 8'b1100111;
DRAM[59883] = 8'b1100111;
DRAM[59884] = 8'b1100111;
DRAM[59885] = 8'b1101000;
DRAM[59886] = 8'b1101001;
DRAM[59887] = 8'b1101010;
DRAM[59888] = 8'b1101101;
DRAM[59889] = 8'b1101100;
DRAM[59890] = 8'b1101100;
DRAM[59891] = 8'b1101101;
DRAM[59892] = 8'b1101111;
DRAM[59893] = 8'b1110001;
DRAM[59894] = 8'b1110000;
DRAM[59895] = 8'b1101111;
DRAM[59896] = 8'b1101100;
DRAM[59897] = 8'b1101100;
DRAM[59898] = 8'b1101100;
DRAM[59899] = 8'b1101011;
DRAM[59900] = 8'b1101010;
DRAM[59901] = 8'b1101001;
DRAM[59902] = 8'b1100111;
DRAM[59903] = 8'b1100110;
DRAM[59904] = 8'b10010110;
DRAM[59905] = 8'b10010100;
DRAM[59906] = 8'b10010001;
DRAM[59907] = 8'b10001111;
DRAM[59908] = 8'b10001110;
DRAM[59909] = 8'b10001111;
DRAM[59910] = 8'b10010000;
DRAM[59911] = 8'b10010001;
DRAM[59912] = 8'b10001001;
DRAM[59913] = 8'b10001110;
DRAM[59914] = 8'b10010100;
DRAM[59915] = 8'b10100001;
DRAM[59916] = 8'b10111100;
DRAM[59917] = 8'b11011110;
DRAM[59918] = 8'b11110010;
DRAM[59919] = 8'b11110111;
DRAM[59920] = 8'b11111011;
DRAM[59921] = 8'b11111100;
DRAM[59922] = 8'b11111101;
DRAM[59923] = 8'b11111101;
DRAM[59924] = 8'b11111011;
DRAM[59925] = 8'b11111000;
DRAM[59926] = 8'b11110100;
DRAM[59927] = 8'b11110010;
DRAM[59928] = 8'b11110011;
DRAM[59929] = 8'b11110000;
DRAM[59930] = 8'b11101100;
DRAM[59931] = 8'b11101010;
DRAM[59932] = 8'b11101011;
DRAM[59933] = 8'b11101100;
DRAM[59934] = 8'b11101100;
DRAM[59935] = 8'b11101100;
DRAM[59936] = 8'b11100110;
DRAM[59937] = 8'b11100100;
DRAM[59938] = 8'b11100000;
DRAM[59939] = 8'b11011110;
DRAM[59940] = 8'b11011100;
DRAM[59941] = 8'b11011010;
DRAM[59942] = 8'b11010110;
DRAM[59943] = 8'b11010100;
DRAM[59944] = 8'b11001101;
DRAM[59945] = 8'b11001100;
DRAM[59946] = 8'b11001010;
DRAM[59947] = 8'b11000111;
DRAM[59948] = 8'b11000011;
DRAM[59949] = 8'b10111111;
DRAM[59950] = 8'b10111100;
DRAM[59951] = 8'b10111001;
DRAM[59952] = 8'b10111001;
DRAM[59953] = 8'b10110100;
DRAM[59954] = 8'b10101111;
DRAM[59955] = 8'b10101101;
DRAM[59956] = 8'b10101101;
DRAM[59957] = 8'b10101010;
DRAM[59958] = 8'b10100010;
DRAM[59959] = 8'b10011100;
DRAM[59960] = 8'b10100101;
DRAM[59961] = 8'b10011001;
DRAM[59962] = 8'b10001101;
DRAM[59963] = 8'b10001110;
DRAM[59964] = 8'b10011011;
DRAM[59965] = 8'b10100010;
DRAM[59966] = 8'b10010110;
DRAM[59967] = 8'b10000100;
DRAM[59968] = 8'b10010011;
DRAM[59969] = 8'b10011001;
DRAM[59970] = 8'b10011111;
DRAM[59971] = 8'b10100010;
DRAM[59972] = 8'b10011110;
DRAM[59973] = 8'b10011001;
DRAM[59974] = 8'b10010101;
DRAM[59975] = 8'b10010100;
DRAM[59976] = 8'b10010101;
DRAM[59977] = 8'b10011011;
DRAM[59978] = 8'b10010101;
DRAM[59979] = 8'b10010000;
DRAM[59980] = 8'b10010111;
DRAM[59981] = 8'b10011000;
DRAM[59982] = 8'b10001100;
DRAM[59983] = 8'b10000010;
DRAM[59984] = 8'b10000111;
DRAM[59985] = 8'b10000101;
DRAM[59986] = 8'b10000000;
DRAM[59987] = 8'b10000010;
DRAM[59988] = 8'b10000011;
DRAM[59989] = 8'b1110111;
DRAM[59990] = 8'b1110011;
DRAM[59991] = 8'b1111101;
DRAM[59992] = 8'b1111110;
DRAM[59993] = 8'b1111100;
DRAM[59994] = 8'b1110111;
DRAM[59995] = 8'b1101011;
DRAM[59996] = 8'b1110001;
DRAM[59997] = 8'b1110110;
DRAM[59998] = 8'b1101000;
DRAM[59999] = 8'b1101011;
DRAM[60000] = 8'b10000001;
DRAM[60001] = 8'b1110011;
DRAM[60002] = 8'b1110111;
DRAM[60003] = 8'b1110100;
DRAM[60004] = 8'b1111000;
DRAM[60005] = 8'b1111110;
DRAM[60006] = 8'b1110110;
DRAM[60007] = 8'b1111110;
DRAM[60008] = 8'b1101000;
DRAM[60009] = 8'b1110101;
DRAM[60010] = 8'b1111110;
DRAM[60011] = 8'b1111011;
DRAM[60012] = 8'b1110100;
DRAM[60013] = 8'b1110011;
DRAM[60014] = 8'b1111000;
DRAM[60015] = 8'b1111101;
DRAM[60016] = 8'b1110011;
DRAM[60017] = 8'b1110101;
DRAM[60018] = 8'b1110110;
DRAM[60019] = 8'b1110111;
DRAM[60020] = 8'b1110111;
DRAM[60021] = 8'b1111000;
DRAM[60022] = 8'b1111011;
DRAM[60023] = 8'b1111101;
DRAM[60024] = 8'b1111110;
DRAM[60025] = 8'b10000101;
DRAM[60026] = 8'b1110100;
DRAM[60027] = 8'b1110110;
DRAM[60028] = 8'b1111100;
DRAM[60029] = 8'b1110000;
DRAM[60030] = 8'b1101111;
DRAM[60031] = 8'b1101010;
DRAM[60032] = 8'b1110001;
DRAM[60033] = 8'b1100110;
DRAM[60034] = 8'b1101111;
DRAM[60035] = 8'b1101110;
DRAM[60036] = 8'b1101110;
DRAM[60037] = 8'b1101111;
DRAM[60038] = 8'b1101010;
DRAM[60039] = 8'b1111000;
DRAM[60040] = 8'b1111010;
DRAM[60041] = 8'b1111001;
DRAM[60042] = 8'b1110001;
DRAM[60043] = 8'b1101001;
DRAM[60044] = 8'b1101011;
DRAM[60045] = 8'b1110101;
DRAM[60046] = 8'b1111000;
DRAM[60047] = 8'b1110100;
DRAM[60048] = 8'b1100011;
DRAM[60049] = 8'b1101100;
DRAM[60050] = 8'b1110100;
DRAM[60051] = 8'b1110110;
DRAM[60052] = 8'b1110100;
DRAM[60053] = 8'b1110010;
DRAM[60054] = 8'b1110100;
DRAM[60055] = 8'b1111010;
DRAM[60056] = 8'b1110011;
DRAM[60057] = 8'b1110011;
DRAM[60058] = 8'b1110000;
DRAM[60059] = 8'b1101110;
DRAM[60060] = 8'b1110110;
DRAM[60061] = 8'b10000001;
DRAM[60062] = 8'b1111111;
DRAM[60063] = 8'b1110110;
DRAM[60064] = 8'b1110101;
DRAM[60065] = 8'b1101111;
DRAM[60066] = 8'b1110111;
DRAM[60067] = 8'b1110001;
DRAM[60068] = 8'b1110000;
DRAM[60069] = 8'b1110100;
DRAM[60070] = 8'b1101010;
DRAM[60071] = 8'b1110000;
DRAM[60072] = 8'b1111101;
DRAM[60073] = 8'b10000000;
DRAM[60074] = 8'b10000001;
DRAM[60075] = 8'b1111110;
DRAM[60076] = 8'b1111001;
DRAM[60077] = 8'b1111011;
DRAM[60078] = 8'b10000100;
DRAM[60079] = 8'b10001100;
DRAM[60080] = 8'b10011010;
DRAM[60081] = 8'b10011011;
DRAM[60082] = 8'b10100000;
DRAM[60083] = 8'b10101000;
DRAM[60084] = 8'b10101110;
DRAM[60085] = 8'b10110010;
DRAM[60086] = 8'b10111010;
DRAM[60087] = 8'b11000010;
DRAM[60088] = 8'b11001000;
DRAM[60089] = 8'b11001110;
DRAM[60090] = 8'b11010101;
DRAM[60091] = 8'b11011100;
DRAM[60092] = 8'b11100001;
DRAM[60093] = 8'b11101001;
DRAM[60094] = 8'b11110001;
DRAM[60095] = 8'b11111000;
DRAM[60096] = 8'b11110111;
DRAM[60097] = 8'b11110100;
DRAM[60098] = 8'b11100000;
DRAM[60099] = 8'b10111100;
DRAM[60100] = 8'b10011101;
DRAM[60101] = 8'b10010010;
DRAM[60102] = 8'b10010001;
DRAM[60103] = 8'b10010000;
DRAM[60104] = 8'b10010011;
DRAM[60105] = 8'b10010011;
DRAM[60106] = 8'b10010001;
DRAM[60107] = 8'b10001111;
DRAM[60108] = 8'b10001100;
DRAM[60109] = 8'b10001000;
DRAM[60110] = 8'b10000101;
DRAM[60111] = 8'b10000100;
DRAM[60112] = 8'b1111111;
DRAM[60113] = 8'b1111101;
DRAM[60114] = 8'b1111001;
DRAM[60115] = 8'b1110110;
DRAM[60116] = 8'b1110100;
DRAM[60117] = 8'b1110100;
DRAM[60118] = 8'b1110100;
DRAM[60119] = 8'b1110101;
DRAM[60120] = 8'b1110111;
DRAM[60121] = 8'b1110110;
DRAM[60122] = 8'b1110101;
DRAM[60123] = 8'b1110011;
DRAM[60124] = 8'b1110010;
DRAM[60125] = 8'b1110000;
DRAM[60126] = 8'b1101111;
DRAM[60127] = 8'b1101111;
DRAM[60128] = 8'b1101011;
DRAM[60129] = 8'b1101011;
DRAM[60130] = 8'b1101010;
DRAM[60131] = 8'b1101001;
DRAM[60132] = 8'b1101001;
DRAM[60133] = 8'b1101001;
DRAM[60134] = 8'b1101001;
DRAM[60135] = 8'b1101001;
DRAM[60136] = 8'b1101000;
DRAM[60137] = 8'b1100111;
DRAM[60138] = 8'b1100111;
DRAM[60139] = 8'b1100111;
DRAM[60140] = 8'b1100111;
DRAM[60141] = 8'b1101000;
DRAM[60142] = 8'b1101001;
DRAM[60143] = 8'b1101010;
DRAM[60144] = 8'b1101100;
DRAM[60145] = 8'b1101100;
DRAM[60146] = 8'b1101100;
DRAM[60147] = 8'b1101110;
DRAM[60148] = 8'b1110000;
DRAM[60149] = 8'b1110001;
DRAM[60150] = 8'b1110000;
DRAM[60151] = 8'b1101110;
DRAM[60152] = 8'b1101100;
DRAM[60153] = 8'b1101100;
DRAM[60154] = 8'b1101100;
DRAM[60155] = 8'b1101011;
DRAM[60156] = 8'b1101010;
DRAM[60157] = 8'b1101001;
DRAM[60158] = 8'b1100111;
DRAM[60159] = 8'b1100110;
DRAM[60160] = 8'b10010101;
DRAM[60161] = 8'b10010011;
DRAM[60162] = 8'b10010000;
DRAM[60163] = 8'b10001110;
DRAM[60164] = 8'b10001100;
DRAM[60165] = 8'b10001101;
DRAM[60166] = 8'b10001111;
DRAM[60167] = 8'b10010000;
DRAM[60168] = 8'b10010001;
DRAM[60169] = 8'b10010011;
DRAM[60170] = 8'b10011000;
DRAM[60171] = 8'b10101000;
DRAM[60172] = 8'b11000100;
DRAM[60173] = 8'b11100010;
DRAM[60174] = 8'b11110001;
DRAM[60175] = 8'b11110010;
DRAM[60176] = 8'b11111011;
DRAM[60177] = 8'b11111011;
DRAM[60178] = 8'b11111011;
DRAM[60179] = 8'b11111011;
DRAM[60180] = 8'b11111010;
DRAM[60181] = 8'b11111000;
DRAM[60182] = 8'b11110100;
DRAM[60183] = 8'b11110010;
DRAM[60184] = 8'b11101110;
DRAM[60185] = 8'b11101100;
DRAM[60186] = 8'b11101010;
DRAM[60187] = 8'b11101011;
DRAM[60188] = 8'b11101101;
DRAM[60189] = 8'b11101110;
DRAM[60190] = 8'b11101110;
DRAM[60191] = 8'b11101101;
DRAM[60192] = 8'b11101011;
DRAM[60193] = 8'b11100101;
DRAM[60194] = 8'b11011011;
DRAM[60195] = 8'b11010101;
DRAM[60196] = 8'b11010011;
DRAM[60197] = 8'b11010110;
DRAM[60198] = 8'b11011000;
DRAM[60199] = 8'b11011010;
DRAM[60200] = 8'b11010000;
DRAM[60201] = 8'b11001110;
DRAM[60202] = 8'b11001011;
DRAM[60203] = 8'b11000111;
DRAM[60204] = 8'b11000010;
DRAM[60205] = 8'b10111101;
DRAM[60206] = 8'b10111010;
DRAM[60207] = 8'b10111000;
DRAM[60208] = 8'b10101001;
DRAM[60209] = 8'b10101000;
DRAM[60210] = 8'b10101001;
DRAM[60211] = 8'b10101100;
DRAM[60212] = 8'b10110000;
DRAM[60213] = 8'b10101110;
DRAM[60214] = 8'b10101000;
DRAM[60215] = 8'b10100001;
DRAM[60216] = 8'b10001101;
DRAM[60217] = 8'b10001110;
DRAM[60218] = 8'b10001100;
DRAM[60219] = 8'b10001000;
DRAM[60220] = 8'b10000100;
DRAM[60221] = 8'b10000010;
DRAM[60222] = 8'b10000010;
DRAM[60223] = 8'b10000001;
DRAM[60224] = 8'b1111110;
DRAM[60225] = 8'b10000110;
DRAM[60226] = 8'b10010000;
DRAM[60227] = 8'b10001111;
DRAM[60228] = 8'b1111111;
DRAM[60229] = 8'b1110100;
DRAM[60230] = 8'b10000000;
DRAM[60231] = 8'b10010100;
DRAM[60232] = 8'b10001101;
DRAM[60233] = 8'b10100011;
DRAM[60234] = 8'b10100001;
DRAM[60235] = 8'b10010110;
DRAM[60236] = 8'b10010110;
DRAM[60237] = 8'b10001101;
DRAM[60238] = 8'b10000010;
DRAM[60239] = 8'b10001011;
DRAM[60240] = 8'b10000111;
DRAM[60241] = 8'b10001101;
DRAM[60242] = 8'b10000100;
DRAM[60243] = 8'b1111111;
DRAM[60244] = 8'b10000110;
DRAM[60245] = 8'b1111011;
DRAM[60246] = 8'b1110011;
DRAM[60247] = 8'b10000100;
DRAM[60248] = 8'b1111100;
DRAM[60249] = 8'b1110101;
DRAM[60250] = 8'b1111011;
DRAM[60251] = 8'b1101000;
DRAM[60252] = 8'b1101101;
DRAM[60253] = 8'b1110110;
DRAM[60254] = 8'b1011101;
DRAM[60255] = 8'b1100101;
DRAM[60256] = 8'b1101011;
DRAM[60257] = 8'b1101011;
DRAM[60258] = 8'b1110111;
DRAM[60259] = 8'b1110010;
DRAM[60260] = 8'b1110111;
DRAM[60261] = 8'b10000011;
DRAM[60262] = 8'b1111000;
DRAM[60263] = 8'b1110111;
DRAM[60264] = 8'b1110101;
DRAM[60265] = 8'b1110011;
DRAM[60266] = 8'b1110010;
DRAM[60267] = 8'b1110011;
DRAM[60268] = 8'b1111000;
DRAM[60269] = 8'b1111010;
DRAM[60270] = 8'b1110111;
DRAM[60271] = 8'b1110010;
DRAM[60272] = 8'b1111101;
DRAM[60273] = 8'b1110111;
DRAM[60274] = 8'b1110001;
DRAM[60275] = 8'b1110011;
DRAM[60276] = 8'b1111001;
DRAM[60277] = 8'b1111110;
DRAM[60278] = 8'b1111110;
DRAM[60279] = 8'b1111011;
DRAM[60280] = 8'b10000001;
DRAM[60281] = 8'b10000010;
DRAM[60282] = 8'b1110001;
DRAM[60283] = 8'b1111001;
DRAM[60284] = 8'b1111111;
DRAM[60285] = 8'b1101110;
DRAM[60286] = 8'b1101011;
DRAM[60287] = 8'b1101010;
DRAM[60288] = 8'b1110001;
DRAM[60289] = 8'b1100010;
DRAM[60290] = 8'b1101011;
DRAM[60291] = 8'b1101110;
DRAM[60292] = 8'b1101111;
DRAM[60293] = 8'b1101101;
DRAM[60294] = 8'b1100110;
DRAM[60295] = 8'b1111000;
DRAM[60296] = 8'b1110110;
DRAM[60297] = 8'b1111000;
DRAM[60298] = 8'b1110010;
DRAM[60299] = 8'b1100111;
DRAM[60300] = 8'b1101001;
DRAM[60301] = 8'b1110100;
DRAM[60302] = 8'b1110111;
DRAM[60303] = 8'b1110001;
DRAM[60304] = 8'b1101110;
DRAM[60305] = 8'b1101101;
DRAM[60306] = 8'b1110100;
DRAM[60307] = 8'b1110111;
DRAM[60308] = 8'b1110000;
DRAM[60309] = 8'b1110000;
DRAM[60310] = 8'b1110101;
DRAM[60311] = 8'b1110010;
DRAM[60312] = 8'b1110011;
DRAM[60313] = 8'b1111000;
DRAM[60314] = 8'b1111000;
DRAM[60315] = 8'b1110011;
DRAM[60316] = 8'b1110100;
DRAM[60317] = 8'b1111011;
DRAM[60318] = 8'b10000000;
DRAM[60319] = 8'b10000000;
DRAM[60320] = 8'b1111001;
DRAM[60321] = 8'b1110011;
DRAM[60322] = 8'b1111101;
DRAM[60323] = 8'b1111000;
DRAM[60324] = 8'b1111000;
DRAM[60325] = 8'b1111100;
DRAM[60326] = 8'b1101111;
DRAM[60327] = 8'b1110010;
DRAM[60328] = 8'b1111001;
DRAM[60329] = 8'b1111101;
DRAM[60330] = 8'b10000001;
DRAM[60331] = 8'b10000010;
DRAM[60332] = 8'b10000001;
DRAM[60333] = 8'b10000011;
DRAM[60334] = 8'b10001001;
DRAM[60335] = 8'b10001110;
DRAM[60336] = 8'b10010011;
DRAM[60337] = 8'b10010011;
DRAM[60338] = 8'b10011010;
DRAM[60339] = 8'b10100100;
DRAM[60340] = 8'b10101100;
DRAM[60341] = 8'b10110100;
DRAM[60342] = 8'b10111110;
DRAM[60343] = 8'b11001000;
DRAM[60344] = 8'b11001011;
DRAM[60345] = 8'b11010010;
DRAM[60346] = 8'b11011001;
DRAM[60347] = 8'b11011110;
DRAM[60348] = 8'b11100000;
DRAM[60349] = 8'b11100110;
DRAM[60350] = 8'b11110000;
DRAM[60351] = 8'b11111000;
DRAM[60352] = 8'b11110100;
DRAM[60353] = 8'b11110101;
DRAM[60354] = 8'b11101000;
DRAM[60355] = 8'b11001010;
DRAM[60356] = 8'b10101011;
DRAM[60357] = 8'b10011001;
DRAM[60358] = 8'b10010001;
DRAM[60359] = 8'b10001110;
DRAM[60360] = 8'b10010100;
DRAM[60361] = 8'b10010011;
DRAM[60362] = 8'b10010010;
DRAM[60363] = 8'b10001111;
DRAM[60364] = 8'b10001100;
DRAM[60365] = 8'b10001001;
DRAM[60366] = 8'b10000110;
DRAM[60367] = 8'b10000100;
DRAM[60368] = 8'b1111111;
DRAM[60369] = 8'b1111100;
DRAM[60370] = 8'b1111000;
DRAM[60371] = 8'b1110100;
DRAM[60372] = 8'b1110010;
DRAM[60373] = 8'b1110010;
DRAM[60374] = 8'b1110100;
DRAM[60375] = 8'b1110101;
DRAM[60376] = 8'b1110110;
DRAM[60377] = 8'b1110101;
DRAM[60378] = 8'b1110101;
DRAM[60379] = 8'b1110011;
DRAM[60380] = 8'b1110010;
DRAM[60381] = 8'b1110001;
DRAM[60382] = 8'b1110000;
DRAM[60383] = 8'b1101111;
DRAM[60384] = 8'b1101011;
DRAM[60385] = 8'b1101010;
DRAM[60386] = 8'b1101001;
DRAM[60387] = 8'b1101001;
DRAM[60388] = 8'b1101000;
DRAM[60389] = 8'b1101000;
DRAM[60390] = 8'b1101001;
DRAM[60391] = 8'b1101001;
DRAM[60392] = 8'b1101000;
DRAM[60393] = 8'b1100111;
DRAM[60394] = 8'b1100111;
DRAM[60395] = 8'b1100111;
DRAM[60396] = 8'b1100111;
DRAM[60397] = 8'b1101000;
DRAM[60398] = 8'b1101001;
DRAM[60399] = 8'b1101010;
DRAM[60400] = 8'b1101100;
DRAM[60401] = 8'b1101011;
DRAM[60402] = 8'b1101100;
DRAM[60403] = 8'b1101110;
DRAM[60404] = 8'b1110001;
DRAM[60405] = 8'b1110001;
DRAM[60406] = 8'b1101111;
DRAM[60407] = 8'b1101110;
DRAM[60408] = 8'b1101100;
DRAM[60409] = 8'b1101100;
DRAM[60410] = 8'b1101100;
DRAM[60411] = 8'b1101011;
DRAM[60412] = 8'b1101010;
DRAM[60413] = 8'b1101001;
DRAM[60414] = 8'b1100111;
DRAM[60415] = 8'b1100110;
DRAM[60416] = 8'b10010110;
DRAM[60417] = 8'b10010100;
DRAM[60418] = 8'b10010001;
DRAM[60419] = 8'b10001111;
DRAM[60420] = 8'b10001101;
DRAM[60421] = 8'b10001101;
DRAM[60422] = 8'b10001110;
DRAM[60423] = 8'b10001111;
DRAM[60424] = 8'b10010100;
DRAM[60425] = 8'b10010101;
DRAM[60426] = 8'b10011100;
DRAM[60427] = 8'b10110000;
DRAM[60428] = 8'b11001110;
DRAM[60429] = 8'b11101000;
DRAM[60430] = 8'b11110100;
DRAM[60431] = 8'b11110100;
DRAM[60432] = 8'b11111010;
DRAM[60433] = 8'b11111001;
DRAM[60434] = 8'b11110111;
DRAM[60435] = 8'b11111000;
DRAM[60436] = 8'b11111010;
DRAM[60437] = 8'b11111001;
DRAM[60438] = 8'b11110110;
DRAM[60439] = 8'b11110011;
DRAM[60440] = 8'b11101100;
DRAM[60441] = 8'b11101100;
DRAM[60442] = 8'b11101101;
DRAM[60443] = 8'b11101111;
DRAM[60444] = 8'b11110001;
DRAM[60445] = 8'b11110000;
DRAM[60446] = 8'b11101100;
DRAM[60447] = 8'b11101001;
DRAM[60448] = 8'b11100010;
DRAM[60449] = 8'b11011011;
DRAM[60450] = 8'b11010010;
DRAM[60451] = 8'b11001100;
DRAM[60452] = 8'b11001010;
DRAM[60453] = 8'b11001101;
DRAM[60454] = 8'b11010000;
DRAM[60455] = 8'b11010001;
DRAM[60456] = 8'b11010001;
DRAM[60457] = 8'b11001111;
DRAM[60458] = 8'b11001100;
DRAM[60459] = 8'b11001000;
DRAM[60460] = 8'b11000100;
DRAM[60461] = 8'b11000000;
DRAM[60462] = 8'b10111101;
DRAM[60463] = 8'b10111100;
DRAM[60464] = 8'b10110110;
DRAM[60465] = 8'b10110110;
DRAM[60466] = 8'b10110110;
DRAM[60467] = 8'b10110111;
DRAM[60468] = 8'b10110111;
DRAM[60469] = 8'b10110001;
DRAM[60470] = 8'b10101001;
DRAM[60471] = 8'b10100010;
DRAM[60472] = 8'b10010110;
DRAM[60473] = 8'b10010111;
DRAM[60474] = 8'b10010110;
DRAM[60475] = 8'b10010000;
DRAM[60476] = 8'b10000110;
DRAM[60477] = 8'b1111111;
DRAM[60478] = 8'b10000000;
DRAM[60479] = 8'b10000100;
DRAM[60480] = 8'b1110100;
DRAM[60481] = 8'b1110110;
DRAM[60482] = 8'b1111101;
DRAM[60483] = 8'b10000011;
DRAM[60484] = 8'b1111101;
DRAM[60485] = 8'b1111010;
DRAM[60486] = 8'b10001010;
DRAM[60487] = 8'b10100000;
DRAM[60488] = 8'b10010110;
DRAM[60489] = 8'b10101001;
DRAM[60490] = 8'b10100110;
DRAM[60491] = 8'b10011011;
DRAM[60492] = 8'b10011001;
DRAM[60493] = 8'b10001110;
DRAM[60494] = 8'b10000101;
DRAM[60495] = 8'b10010001;
DRAM[60496] = 8'b1111110;
DRAM[60497] = 8'b10001101;
DRAM[60498] = 8'b10000100;
DRAM[60499] = 8'b1111011;
DRAM[60500] = 8'b10000101;
DRAM[60501] = 8'b10000111;
DRAM[60502] = 8'b10000010;
DRAM[60503] = 8'b10001010;
DRAM[60504] = 8'b1111011;
DRAM[60505] = 8'b1110111;
DRAM[60506] = 8'b1111110;
DRAM[60507] = 8'b1101010;
DRAM[60508] = 8'b1101100;
DRAM[60509] = 8'b1110101;
DRAM[60510] = 8'b1100001;
DRAM[60511] = 8'b1101110;
DRAM[60512] = 8'b1011111;
DRAM[60513] = 8'b1101100;
DRAM[60514] = 8'b1111011;
DRAM[60515] = 8'b1101101;
DRAM[60516] = 8'b1110010;
DRAM[60517] = 8'b10000110;
DRAM[60518] = 8'b1111011;
DRAM[60519] = 8'b1101111;
DRAM[60520] = 8'b1111001;
DRAM[60521] = 8'b1110010;
DRAM[60522] = 8'b1101100;
DRAM[60523] = 8'b1101100;
DRAM[60524] = 8'b1101110;
DRAM[60525] = 8'b1101111;
DRAM[60526] = 8'b1101101;
DRAM[60527] = 8'b1101011;
DRAM[60528] = 8'b1100011;
DRAM[60529] = 8'b1110001;
DRAM[60530] = 8'b10000000;
DRAM[60531] = 8'b10000100;
DRAM[60532] = 8'b1111111;
DRAM[60533] = 8'b1111010;
DRAM[60534] = 8'b1111011;
DRAM[60535] = 8'b1111111;
DRAM[60536] = 8'b1111101;
DRAM[60537] = 8'b1111101;
DRAM[60538] = 8'b1101101;
DRAM[60539] = 8'b1111001;
DRAM[60540] = 8'b10000001;
DRAM[60541] = 8'b1101111;
DRAM[60542] = 8'b1101010;
DRAM[60543] = 8'b1101001;
DRAM[60544] = 8'b1110001;
DRAM[60545] = 8'b1100001;
DRAM[60546] = 8'b1101010;
DRAM[60547] = 8'b1101111;
DRAM[60548] = 8'b1110001;
DRAM[60549] = 8'b1101111;
DRAM[60550] = 8'b1100111;
DRAM[60551] = 8'b1110111;
DRAM[60552] = 8'b1110010;
DRAM[60553] = 8'b1110101;
DRAM[60554] = 8'b1110010;
DRAM[60555] = 8'b1101011;
DRAM[60556] = 8'b1101100;
DRAM[60557] = 8'b1110011;
DRAM[60558] = 8'b1110100;
DRAM[60559] = 8'b1101110;
DRAM[60560] = 8'b1110110;
DRAM[60561] = 8'b1101101;
DRAM[60562] = 8'b1101110;
DRAM[60563] = 8'b1110000;
DRAM[60564] = 8'b1101110;
DRAM[60565] = 8'b1110010;
DRAM[60566] = 8'b1110110;
DRAM[60567] = 8'b1101111;
DRAM[60568] = 8'b10000001;
DRAM[60569] = 8'b1110111;
DRAM[60570] = 8'b1101101;
DRAM[60571] = 8'b1101101;
DRAM[60572] = 8'b1111001;
DRAM[60573] = 8'b10000011;
DRAM[60574] = 8'b1111110;
DRAM[60575] = 8'b1110101;
DRAM[60576] = 8'b1110100;
DRAM[60577] = 8'b1101111;
DRAM[60578] = 8'b1111010;
DRAM[60579] = 8'b1111000;
DRAM[60580] = 8'b1111011;
DRAM[60581] = 8'b10000000;
DRAM[60582] = 8'b1110011;
DRAM[60583] = 8'b1110101;
DRAM[60584] = 8'b10000101;
DRAM[60585] = 8'b10000110;
DRAM[60586] = 8'b10001000;
DRAM[60587] = 8'b10001011;
DRAM[60588] = 8'b10001100;
DRAM[60589] = 8'b10001011;
DRAM[60590] = 8'b10001000;
DRAM[60591] = 8'b10000110;
DRAM[60592] = 8'b10010010;
DRAM[60593] = 8'b10010011;
DRAM[60594] = 8'b10011001;
DRAM[60595] = 8'b10100011;
DRAM[60596] = 8'b10101100;
DRAM[60597] = 8'b10110011;
DRAM[60598] = 8'b10111101;
DRAM[60599] = 8'b11000111;
DRAM[60600] = 8'b11001111;
DRAM[60601] = 8'b11010101;
DRAM[60602] = 8'b11011101;
DRAM[60603] = 8'b11100001;
DRAM[60604] = 8'b11100010;
DRAM[60605] = 8'b11100111;
DRAM[60606] = 8'b11101111;
DRAM[60607] = 8'b11110111;
DRAM[60608] = 8'b11110110;
DRAM[60609] = 8'b11110111;
DRAM[60610] = 8'b11101101;
DRAM[60611] = 8'b11010100;
DRAM[60612] = 8'b10110111;
DRAM[60613] = 8'b10100011;
DRAM[60614] = 8'b10011010;
DRAM[60615] = 8'b10010110;
DRAM[60616] = 8'b10010011;
DRAM[60617] = 8'b10010011;
DRAM[60618] = 8'b10010001;
DRAM[60619] = 8'b10001111;
DRAM[60620] = 8'b10001101;
DRAM[60621] = 8'b10001010;
DRAM[60622] = 8'b10000111;
DRAM[60623] = 8'b10000110;
DRAM[60624] = 8'b10000000;
DRAM[60625] = 8'b1111101;
DRAM[60626] = 8'b1111001;
DRAM[60627] = 8'b1110101;
DRAM[60628] = 8'b1110011;
DRAM[60629] = 8'b1110011;
DRAM[60630] = 8'b1110100;
DRAM[60631] = 8'b1110101;
DRAM[60632] = 8'b1110101;
DRAM[60633] = 8'b1110100;
DRAM[60634] = 8'b1110011;
DRAM[60635] = 8'b1110010;
DRAM[60636] = 8'b1110001;
DRAM[60637] = 8'b1110000;
DRAM[60638] = 8'b1101111;
DRAM[60639] = 8'b1101111;
DRAM[60640] = 8'b1101011;
DRAM[60641] = 8'b1101010;
DRAM[60642] = 8'b1101001;
DRAM[60643] = 8'b1101000;
DRAM[60644] = 8'b1101000;
DRAM[60645] = 8'b1101000;
DRAM[60646] = 8'b1101000;
DRAM[60647] = 8'b1101001;
DRAM[60648] = 8'b1101000;
DRAM[60649] = 8'b1100111;
DRAM[60650] = 8'b1100111;
DRAM[60651] = 8'b1100111;
DRAM[60652] = 8'b1100111;
DRAM[60653] = 8'b1101000;
DRAM[60654] = 8'b1101001;
DRAM[60655] = 8'b1101010;
DRAM[60656] = 8'b1101011;
DRAM[60657] = 8'b1101011;
DRAM[60658] = 8'b1101100;
DRAM[60659] = 8'b1101111;
DRAM[60660] = 8'b1110001;
DRAM[60661] = 8'b1110001;
DRAM[60662] = 8'b1101111;
DRAM[60663] = 8'b1101101;
DRAM[60664] = 8'b1101100;
DRAM[60665] = 8'b1101100;
DRAM[60666] = 8'b1101100;
DRAM[60667] = 8'b1101011;
DRAM[60668] = 8'b1101010;
DRAM[60669] = 8'b1101001;
DRAM[60670] = 8'b1100111;
DRAM[60671] = 8'b1100110;
DRAM[60672] = 8'b10010111;
DRAM[60673] = 8'b10010110;
DRAM[60674] = 8'b10010100;
DRAM[60675] = 8'b10010010;
DRAM[60676] = 8'b10010001;
DRAM[60677] = 8'b10010000;
DRAM[60678] = 8'b10001111;
DRAM[60679] = 8'b10001111;
DRAM[60680] = 8'b10010001;
DRAM[60681] = 8'b10010011;
DRAM[60682] = 8'b10011111;
DRAM[60683] = 8'b10110111;
DRAM[60684] = 8'b11010101;
DRAM[60685] = 8'b11101110;
DRAM[60686] = 8'b11111001;
DRAM[60687] = 8'b11111010;
DRAM[60688] = 8'b11111010;
DRAM[60689] = 8'b11110111;
DRAM[60690] = 8'b11110101;
DRAM[60691] = 8'b11110110;
DRAM[60692] = 8'b11111001;
DRAM[60693] = 8'b11111001;
DRAM[60694] = 8'b11110110;
DRAM[60695] = 8'b11110010;
DRAM[60696] = 8'b11110000;
DRAM[60697] = 8'b11110000;
DRAM[60698] = 8'b11110001;
DRAM[60699] = 8'b11110010;
DRAM[60700] = 8'b11110001;
DRAM[60701] = 8'b11101101;
DRAM[60702] = 8'b11100110;
DRAM[60703] = 8'b11100010;
DRAM[60704] = 8'b11011101;
DRAM[60705] = 8'b11011011;
DRAM[60706] = 8'b11011000;
DRAM[60707] = 8'b11010110;
DRAM[60708] = 8'b11010101;
DRAM[60709] = 8'b11010011;
DRAM[60710] = 8'b11010000;
DRAM[60711] = 8'b11001110;
DRAM[60712] = 8'b11001100;
DRAM[60713] = 8'b11001010;
DRAM[60714] = 8'b11001000;
DRAM[60715] = 8'b11000110;
DRAM[60716] = 8'b11000100;
DRAM[60717] = 8'b11000010;
DRAM[60718] = 8'b11000010;
DRAM[60719] = 8'b11000010;
DRAM[60720] = 8'b11000110;
DRAM[60721] = 8'b11000101;
DRAM[60722] = 8'b11000100;
DRAM[60723] = 8'b11000011;
DRAM[60724] = 8'b11000000;
DRAM[60725] = 8'b10111001;
DRAM[60726] = 8'b10110000;
DRAM[60727] = 8'b10101001;
DRAM[60728] = 8'b10110001;
DRAM[60729] = 8'b10100001;
DRAM[60730] = 8'b10010100;
DRAM[60731] = 8'b10010011;
DRAM[60732] = 8'b10010110;
DRAM[60733] = 8'b10010010;
DRAM[60734] = 8'b10000111;
DRAM[60735] = 8'b1111110;
DRAM[60736] = 8'b10000001;
DRAM[60737] = 8'b1110111;
DRAM[60738] = 8'b1110101;
DRAM[60739] = 8'b10000000;
DRAM[60740] = 8'b10001011;
DRAM[60741] = 8'b10001110;
DRAM[60742] = 8'b10010000;
DRAM[60743] = 8'b10010011;
DRAM[60744] = 8'b10011101;
DRAM[60745] = 8'b10011111;
DRAM[60746] = 8'b10011010;
DRAM[60747] = 8'b10010110;
DRAM[60748] = 8'b10011001;
DRAM[60749] = 8'b10010100;
DRAM[60750] = 8'b10001010;
DRAM[60751] = 8'b10001001;
DRAM[60752] = 8'b10000110;
DRAM[60753] = 8'b10001110;
DRAM[60754] = 8'b10000111;
DRAM[60755] = 8'b1111101;
DRAM[60756] = 8'b10000001;
DRAM[60757] = 8'b10000110;
DRAM[60758] = 8'b10000010;
DRAM[60759] = 8'b1111110;
DRAM[60760] = 8'b1111110;
DRAM[60761] = 8'b10000000;
DRAM[60762] = 8'b1111110;
DRAM[60763] = 8'b1110000;
DRAM[60764] = 8'b1110011;
DRAM[60765] = 8'b1110111;
DRAM[60766] = 8'b1101111;
DRAM[60767] = 8'b1111000;
DRAM[60768] = 8'b1101001;
DRAM[60769] = 8'b1110011;
DRAM[60770] = 8'b1111100;
DRAM[60771] = 8'b1101001;
DRAM[60772] = 8'b1101011;
DRAM[60773] = 8'b10000001;
DRAM[60774] = 8'b1111010;
DRAM[60775] = 8'b1110010;
DRAM[60776] = 8'b1110110;
DRAM[60777] = 8'b1110111;
DRAM[60778] = 8'b1111000;
DRAM[60779] = 8'b1110001;
DRAM[60780] = 8'b1100101;
DRAM[60781] = 8'b1011110;
DRAM[60782] = 8'b1100110;
DRAM[60783] = 8'b1110010;
DRAM[60784] = 8'b1100101;
DRAM[60785] = 8'b1101011;
DRAM[60786] = 8'b1110011;
DRAM[60787] = 8'b1111010;
DRAM[60788] = 8'b1111110;
DRAM[60789] = 8'b10000001;
DRAM[60790] = 8'b10000011;
DRAM[60791] = 8'b10000101;
DRAM[60792] = 8'b1111001;
DRAM[60793] = 8'b1111011;
DRAM[60794] = 8'b1101011;
DRAM[60795] = 8'b1110111;
DRAM[60796] = 8'b10000001;
DRAM[60797] = 8'b1110010;
DRAM[60798] = 8'b1101101;
DRAM[60799] = 8'b1101001;
DRAM[60800] = 8'b1110001;
DRAM[60801] = 8'b1100101;
DRAM[60802] = 8'b1101110;
DRAM[60803] = 8'b1101111;
DRAM[60804] = 8'b1110010;
DRAM[60805] = 8'b1110101;
DRAM[60806] = 8'b1101100;
DRAM[60807] = 8'b1110111;
DRAM[60808] = 8'b1110011;
DRAM[60809] = 8'b1110011;
DRAM[60810] = 8'b1110011;
DRAM[60811] = 8'b1110010;
DRAM[60812] = 8'b1110010;
DRAM[60813] = 8'b1110010;
DRAM[60814] = 8'b1110001;
DRAM[60815] = 8'b1110001;
DRAM[60816] = 8'b1110011;
DRAM[60817] = 8'b1101110;
DRAM[60818] = 8'b1100111;
DRAM[60819] = 8'b1101000;
DRAM[60820] = 8'b1110000;
DRAM[60821] = 8'b1110101;
DRAM[60822] = 8'b1110100;
DRAM[60823] = 8'b1110010;
DRAM[60824] = 8'b1111011;
DRAM[60825] = 8'b1110110;
DRAM[60826] = 8'b1110001;
DRAM[60827] = 8'b1110000;
DRAM[60828] = 8'b1110011;
DRAM[60829] = 8'b1110110;
DRAM[60830] = 8'b1110111;
DRAM[60831] = 8'b1110101;
DRAM[60832] = 8'b1110101;
DRAM[60833] = 8'b1101101;
DRAM[60834] = 8'b1110110;
DRAM[60835] = 8'b1110011;
DRAM[60836] = 8'b1111001;
DRAM[60837] = 8'b10000010;
DRAM[60838] = 8'b1111001;
DRAM[60839] = 8'b1111101;
DRAM[60840] = 8'b10000111;
DRAM[60841] = 8'b10001000;
DRAM[60842] = 8'b10001011;
DRAM[60843] = 8'b10001111;
DRAM[60844] = 8'b10010011;
DRAM[60845] = 8'b10010011;
DRAM[60846] = 8'b10001111;
DRAM[60847] = 8'b10001010;
DRAM[60848] = 8'b10011000;
DRAM[60849] = 8'b10011000;
DRAM[60850] = 8'b10011110;
DRAM[60851] = 8'b10100110;
DRAM[60852] = 8'b10101100;
DRAM[60853] = 8'b10110000;
DRAM[60854] = 8'b10111000;
DRAM[60855] = 8'b11000000;
DRAM[60856] = 8'b11001101;
DRAM[60857] = 8'b11010011;
DRAM[60858] = 8'b11011011;
DRAM[60859] = 8'b11100001;
DRAM[60860] = 8'b11100101;
DRAM[60861] = 8'b11101001;
DRAM[60862] = 8'b11101111;
DRAM[60863] = 8'b11110100;
DRAM[60864] = 8'b11110110;
DRAM[60865] = 8'b11101111;
DRAM[60866] = 8'b11011111;
DRAM[60867] = 8'b11000111;
DRAM[60868] = 8'b10101111;
DRAM[60869] = 8'b10011111;
DRAM[60870] = 8'b10011010;
DRAM[60871] = 8'b10011010;
DRAM[60872] = 8'b10010100;
DRAM[60873] = 8'b10010011;
DRAM[60874] = 8'b10010010;
DRAM[60875] = 8'b10010000;
DRAM[60876] = 8'b10001101;
DRAM[60877] = 8'b10001010;
DRAM[60878] = 8'b10001000;
DRAM[60879] = 8'b10000110;
DRAM[60880] = 8'b1111111;
DRAM[60881] = 8'b1111101;
DRAM[60882] = 8'b1111010;
DRAM[60883] = 8'b1110110;
DRAM[60884] = 8'b1110100;
DRAM[60885] = 8'b1110100;
DRAM[60886] = 8'b1110100;
DRAM[60887] = 8'b1110101;
DRAM[60888] = 8'b1110011;
DRAM[60889] = 8'b1110010;
DRAM[60890] = 8'b1110010;
DRAM[60891] = 8'b1110001;
DRAM[60892] = 8'b1110000;
DRAM[60893] = 8'b1101111;
DRAM[60894] = 8'b1101110;
DRAM[60895] = 8'b1101110;
DRAM[60896] = 8'b1101010;
DRAM[60897] = 8'b1101010;
DRAM[60898] = 8'b1101001;
DRAM[60899] = 8'b1101000;
DRAM[60900] = 8'b1100111;
DRAM[60901] = 8'b1100111;
DRAM[60902] = 8'b1101000;
DRAM[60903] = 8'b1101000;
DRAM[60904] = 8'b1101000;
DRAM[60905] = 8'b1100111;
DRAM[60906] = 8'b1100111;
DRAM[60907] = 8'b1100111;
DRAM[60908] = 8'b1100111;
DRAM[60909] = 8'b1101000;
DRAM[60910] = 8'b1101001;
DRAM[60911] = 8'b1101010;
DRAM[60912] = 8'b1101011;
DRAM[60913] = 8'b1101011;
DRAM[60914] = 8'b1101100;
DRAM[60915] = 8'b1101111;
DRAM[60916] = 8'b1110010;
DRAM[60917] = 8'b1110010;
DRAM[60918] = 8'b1101111;
DRAM[60919] = 8'b1101100;
DRAM[60920] = 8'b1101100;
DRAM[60921] = 8'b1101100;
DRAM[60922] = 8'b1101100;
DRAM[60923] = 8'b1101011;
DRAM[60924] = 8'b1101010;
DRAM[60925] = 8'b1101001;
DRAM[60926] = 8'b1100111;
DRAM[60927] = 8'b1100110;
DRAM[60928] = 8'b10010101;
DRAM[60929] = 8'b10010101;
DRAM[60930] = 8'b10010100;
DRAM[60931] = 8'b10010100;
DRAM[60932] = 8'b10010010;
DRAM[60933] = 8'b10010000;
DRAM[60934] = 8'b10001101;
DRAM[60935] = 8'b10001100;
DRAM[60936] = 8'b10001111;
DRAM[60937] = 8'b10010100;
DRAM[60938] = 8'b10100010;
DRAM[60939] = 8'b10111100;
DRAM[60940] = 8'b11011001;
DRAM[60941] = 8'b11101110;
DRAM[60942] = 8'b11111000;
DRAM[60943] = 8'b11111011;
DRAM[60944] = 8'b11111101;
DRAM[60945] = 8'b11111001;
DRAM[60946] = 8'b11110101;
DRAM[60947] = 8'b11110101;
DRAM[60948] = 8'b11111000;
DRAM[60949] = 8'b11111000;
DRAM[60950] = 8'b11110100;
DRAM[60951] = 8'b11101111;
DRAM[60952] = 8'b11110010;
DRAM[60953] = 8'b11110001;
DRAM[60954] = 8'b11110000;
DRAM[60955] = 8'b11101111;
DRAM[60956] = 8'b11101101;
DRAM[60957] = 8'b11101001;
DRAM[60958] = 8'b11100100;
DRAM[60959] = 8'b11011111;
DRAM[60960] = 8'b11011111;
DRAM[60961] = 8'b11011101;
DRAM[60962] = 8'b11011011;
DRAM[60963] = 8'b11011011;
DRAM[60964] = 8'b11011010;
DRAM[60965] = 8'b11010111;
DRAM[60966] = 8'b11010011;
DRAM[60967] = 8'b11010000;
DRAM[60968] = 8'b11000110;
DRAM[60969] = 8'b11000101;
DRAM[60970] = 8'b11000011;
DRAM[60971] = 8'b11000001;
DRAM[60972] = 8'b10111111;
DRAM[60973] = 8'b10111111;
DRAM[60974] = 8'b10111111;
DRAM[60975] = 8'b10111111;
DRAM[60976] = 8'b10110110;
DRAM[60977] = 8'b10110110;
DRAM[60978] = 8'b10110101;
DRAM[60979] = 8'b10110100;
DRAM[60980] = 8'b10110010;
DRAM[60981] = 8'b10101110;
DRAM[60982] = 8'b10101001;
DRAM[60983] = 8'b10100101;
DRAM[60984] = 8'b10011000;
DRAM[60985] = 8'b10011000;
DRAM[60986] = 8'b10011000;
DRAM[60987] = 8'b10010001;
DRAM[60988] = 8'b10000011;
DRAM[60989] = 8'b1111000;
DRAM[60990] = 8'b1111011;
DRAM[60991] = 8'b10000101;
DRAM[60992] = 8'b10000010;
DRAM[60993] = 8'b1111001;
DRAM[60994] = 8'b1110010;
DRAM[60995] = 8'b1110101;
DRAM[60996] = 8'b1111101;
DRAM[60997] = 8'b10000001;
DRAM[60998] = 8'b1111110;
DRAM[60999] = 8'b1111010;
DRAM[61000] = 8'b10010011;
DRAM[61001] = 8'b10001110;
DRAM[61002] = 8'b10010011;
DRAM[61003] = 8'b10010111;
DRAM[61004] = 8'b10010010;
DRAM[61005] = 8'b10010000;
DRAM[61006] = 8'b10001110;
DRAM[61007] = 8'b10000110;
DRAM[61008] = 8'b10010110;
DRAM[61009] = 8'b10001001;
DRAM[61010] = 8'b10000101;
DRAM[61011] = 8'b10000111;
DRAM[61012] = 8'b10000011;
DRAM[61013] = 8'b10000001;
DRAM[61014] = 8'b1111110;
DRAM[61015] = 8'b1110110;
DRAM[61016] = 8'b10000000;
DRAM[61017] = 8'b10000111;
DRAM[61018] = 8'b1110111;
DRAM[61019] = 8'b1110100;
DRAM[61020] = 8'b1111011;
DRAM[61021] = 8'b1111001;
DRAM[61022] = 8'b1111011;
DRAM[61023] = 8'b1110111;
DRAM[61024] = 8'b1110011;
DRAM[61025] = 8'b1101111;
DRAM[61026] = 8'b1110111;
DRAM[61027] = 8'b1101110;
DRAM[61028] = 8'b1101110;
DRAM[61029] = 8'b1111000;
DRAM[61030] = 8'b1110011;
DRAM[61031] = 8'b1111001;
DRAM[61032] = 8'b1110101;
DRAM[61033] = 8'b1111001;
DRAM[61034] = 8'b1111100;
DRAM[61035] = 8'b1110110;
DRAM[61036] = 8'b1100110;
DRAM[61037] = 8'b1011100;
DRAM[61038] = 8'b1100011;
DRAM[61039] = 8'b1110010;
DRAM[61040] = 8'b1110100;
DRAM[61041] = 8'b1101011;
DRAM[61042] = 8'b1100100;
DRAM[61043] = 8'b1101010;
DRAM[61044] = 8'b1111010;
DRAM[61045] = 8'b10000101;
DRAM[61046] = 8'b10000111;
DRAM[61047] = 8'b10000011;
DRAM[61048] = 8'b1111010;
DRAM[61049] = 8'b1111110;
DRAM[61050] = 8'b1101100;
DRAM[61051] = 8'b1110011;
DRAM[61052] = 8'b1111110;
DRAM[61053] = 8'b1110101;
DRAM[61054] = 8'b1110010;
DRAM[61055] = 8'b1101010;
DRAM[61056] = 8'b1101111;
DRAM[61057] = 8'b1100111;
DRAM[61058] = 8'b1110000;
DRAM[61059] = 8'b1101101;
DRAM[61060] = 8'b1110001;
DRAM[61061] = 8'b1111001;
DRAM[61062] = 8'b1101111;
DRAM[61063] = 8'b1110100;
DRAM[61064] = 8'b1110110;
DRAM[61065] = 8'b1110000;
DRAM[61066] = 8'b1110000;
DRAM[61067] = 8'b1110110;
DRAM[61068] = 8'b1110101;
DRAM[61069] = 8'b1101110;
DRAM[61070] = 8'b1101110;
DRAM[61071] = 8'b1110101;
DRAM[61072] = 8'b1101100;
DRAM[61073] = 8'b1110010;
DRAM[61074] = 8'b1101000;
DRAM[61075] = 8'b1100101;
DRAM[61076] = 8'b1110011;
DRAM[61077] = 8'b1110010;
DRAM[61078] = 8'b1101011;
DRAM[61079] = 8'b1110011;
DRAM[61080] = 8'b1110000;
DRAM[61081] = 8'b1110110;
DRAM[61082] = 8'b1111010;
DRAM[61083] = 8'b1110110;
DRAM[61084] = 8'b1101101;
DRAM[61085] = 8'b1101010;
DRAM[61086] = 8'b1110010;
DRAM[61087] = 8'b1111100;
DRAM[61088] = 8'b10000010;
DRAM[61089] = 8'b1110101;
DRAM[61090] = 8'b1110110;
DRAM[61091] = 8'b1101111;
DRAM[61092] = 8'b1110101;
DRAM[61093] = 8'b10000011;
DRAM[61094] = 8'b1111111;
DRAM[61095] = 8'b10000111;
DRAM[61096] = 8'b10000011;
DRAM[61097] = 8'b10000110;
DRAM[61098] = 8'b10001100;
DRAM[61099] = 8'b10010001;
DRAM[61100] = 8'b10010110;
DRAM[61101] = 8'b10011001;
DRAM[61102] = 8'b10011100;
DRAM[61103] = 8'b10011110;
DRAM[61104] = 8'b10011100;
DRAM[61105] = 8'b10011100;
DRAM[61106] = 8'b10100010;
DRAM[61107] = 8'b10101001;
DRAM[61108] = 8'b10101110;
DRAM[61109] = 8'b10110000;
DRAM[61110] = 8'b10110101;
DRAM[61111] = 8'b10111100;
DRAM[61112] = 8'b11000101;
DRAM[61113] = 8'b11001011;
DRAM[61114] = 8'b11010011;
DRAM[61115] = 8'b11011101;
DRAM[61116] = 8'b11100101;
DRAM[61117] = 8'b11101011;
DRAM[61118] = 8'b11101111;
DRAM[61119] = 8'b11110001;
DRAM[61120] = 8'b11110100;
DRAM[61121] = 8'b11100111;
DRAM[61122] = 8'b11010011;
DRAM[61123] = 8'b10111100;
DRAM[61124] = 8'b10101000;
DRAM[61125] = 8'b10011010;
DRAM[61126] = 8'b10010110;
DRAM[61127] = 8'b10010110;
DRAM[61128] = 8'b10010110;
DRAM[61129] = 8'b10010101;
DRAM[61130] = 8'b10010011;
DRAM[61131] = 8'b10010001;
DRAM[61132] = 8'b10001101;
DRAM[61133] = 8'b10001001;
DRAM[61134] = 8'b10000110;
DRAM[61135] = 8'b10000100;
DRAM[61136] = 8'b1111101;
DRAM[61137] = 8'b1111100;
DRAM[61138] = 8'b1111001;
DRAM[61139] = 8'b1110111;
DRAM[61140] = 8'b1110101;
DRAM[61141] = 8'b1110100;
DRAM[61142] = 8'b1110011;
DRAM[61143] = 8'b1110011;
DRAM[61144] = 8'b1110001;
DRAM[61145] = 8'b1110000;
DRAM[61146] = 8'b1110000;
DRAM[61147] = 8'b1101111;
DRAM[61148] = 8'b1101110;
DRAM[61149] = 8'b1101110;
DRAM[61150] = 8'b1101101;
DRAM[61151] = 8'b1101101;
DRAM[61152] = 8'b1101010;
DRAM[61153] = 8'b1101001;
DRAM[61154] = 8'b1101000;
DRAM[61155] = 8'b1101000;
DRAM[61156] = 8'b1100111;
DRAM[61157] = 8'b1100111;
DRAM[61158] = 8'b1101000;
DRAM[61159] = 8'b1101000;
DRAM[61160] = 8'b1101000;
DRAM[61161] = 8'b1100111;
DRAM[61162] = 8'b1100111;
DRAM[61163] = 8'b1100111;
DRAM[61164] = 8'b1100111;
DRAM[61165] = 8'b1101000;
DRAM[61166] = 8'b1101001;
DRAM[61167] = 8'b1101010;
DRAM[61168] = 8'b1101010;
DRAM[61169] = 8'b1101011;
DRAM[61170] = 8'b1101101;
DRAM[61171] = 8'b1110000;
DRAM[61172] = 8'b1110010;
DRAM[61173] = 8'b1110010;
DRAM[61174] = 8'b1101111;
DRAM[61175] = 8'b1101100;
DRAM[61176] = 8'b1101100;
DRAM[61177] = 8'b1101100;
DRAM[61178] = 8'b1101100;
DRAM[61179] = 8'b1101011;
DRAM[61180] = 8'b1101010;
DRAM[61181] = 8'b1101001;
DRAM[61182] = 8'b1100111;
DRAM[61183] = 8'b1100110;
DRAM[61184] = 8'b10010001;
DRAM[61185] = 8'b10010010;
DRAM[61186] = 8'b10010010;
DRAM[61187] = 8'b10010010;
DRAM[61188] = 8'b10010000;
DRAM[61189] = 8'b10001101;
DRAM[61190] = 8'b10001010;
DRAM[61191] = 8'b10001000;
DRAM[61192] = 8'b10010001;
DRAM[61193] = 8'b10010110;
DRAM[61194] = 8'b10100110;
DRAM[61195] = 8'b10111111;
DRAM[61196] = 8'b11011001;
DRAM[61197] = 8'b11101011;
DRAM[61198] = 8'b11110100;
DRAM[61199] = 8'b11110111;
DRAM[61200] = 8'b11111111;
DRAM[61201] = 8'b11111011;
DRAM[61202] = 8'b11110110;
DRAM[61203] = 8'b11110101;
DRAM[61204] = 8'b11110111;
DRAM[61205] = 8'b11110110;
DRAM[61206] = 8'b11110001;
DRAM[61207] = 8'b11101100;
DRAM[61208] = 8'b11110000;
DRAM[61209] = 8'b11101110;
DRAM[61210] = 8'b11101100;
DRAM[61211] = 8'b11101011;
DRAM[61212] = 8'b11101010;
DRAM[61213] = 8'b11101000;
DRAM[61214] = 8'b11100101;
DRAM[61215] = 8'b11100011;
DRAM[61216] = 8'b11011010;
DRAM[61217] = 8'b11010110;
DRAM[61218] = 8'b11010000;
DRAM[61219] = 8'b11001100;
DRAM[61220] = 8'b11001011;
DRAM[61221] = 8'b11001100;
DRAM[61222] = 8'b11001100;
DRAM[61223] = 8'b11001100;
DRAM[61224] = 8'b11000101;
DRAM[61225] = 8'b11000011;
DRAM[61226] = 8'b11000000;
DRAM[61227] = 8'b10111101;
DRAM[61228] = 8'b10111010;
DRAM[61229] = 8'b10111000;
DRAM[61230] = 8'b10110111;
DRAM[61231] = 8'b10110111;
DRAM[61232] = 8'b10110100;
DRAM[61233] = 8'b10110100;
DRAM[61234] = 8'b10110011;
DRAM[61235] = 8'b10110001;
DRAM[61236] = 8'b10101111;
DRAM[61237] = 8'b10101011;
DRAM[61238] = 8'b10101000;
DRAM[61239] = 8'b10100110;
DRAM[61240] = 8'b10100111;
DRAM[61241] = 8'b10010100;
DRAM[61242] = 8'b10000111;
DRAM[61243] = 8'b10001100;
DRAM[61244] = 8'b10010101;
DRAM[61245] = 8'b10010011;
DRAM[61246] = 8'b10001010;
DRAM[61247] = 8'b10000011;
DRAM[61248] = 8'b10000110;
DRAM[61249] = 8'b10000111;
DRAM[61250] = 8'b10000100;
DRAM[61251] = 8'b1111100;
DRAM[61252] = 8'b1111000;
DRAM[61253] = 8'b1111101;
DRAM[61254] = 8'b10000111;
DRAM[61255] = 8'b10001101;
DRAM[61256] = 8'b10000110;
DRAM[61257] = 8'b10000111;
DRAM[61258] = 8'b10011100;
DRAM[61259] = 8'b10100010;
DRAM[61260] = 8'b10001110;
DRAM[61261] = 8'b10001010;
DRAM[61262] = 8'b10010100;
DRAM[61263] = 8'b10010001;
DRAM[61264] = 8'b10010111;
DRAM[61265] = 8'b1111010;
DRAM[61266] = 8'b1111100;
DRAM[61267] = 8'b10001111;
DRAM[61268] = 8'b10001010;
DRAM[61269] = 8'b10000100;
DRAM[61270] = 8'b10000110;
DRAM[61271] = 8'b10000001;
DRAM[61272] = 8'b10000000;
DRAM[61273] = 8'b10001010;
DRAM[61274] = 8'b1101110;
DRAM[61275] = 8'b1110100;
DRAM[61276] = 8'b10000000;
DRAM[61277] = 8'b1111001;
DRAM[61278] = 8'b1111111;
DRAM[61279] = 8'b1110001;
DRAM[61280] = 8'b1110011;
DRAM[61281] = 8'b1100100;
DRAM[61282] = 8'b1101111;
DRAM[61283] = 8'b1110110;
DRAM[61284] = 8'b1110111;
DRAM[61285] = 8'b1110011;
DRAM[61286] = 8'b1101011;
DRAM[61287] = 8'b1111110;
DRAM[61288] = 8'b1110110;
DRAM[61289] = 8'b1110001;
DRAM[61290] = 8'b1110000;
DRAM[61291] = 8'b1110000;
DRAM[61292] = 8'b1101001;
DRAM[61293] = 8'b1100000;
DRAM[61294] = 8'b1011111;
DRAM[61295] = 8'b1100101;
DRAM[61296] = 8'b1100101;
DRAM[61297] = 8'b1101101;
DRAM[61298] = 8'b1110110;
DRAM[61299] = 8'b1111010;
DRAM[61300] = 8'b1111010;
DRAM[61301] = 8'b1111001;
DRAM[61302] = 8'b1111011;
DRAM[61303] = 8'b1111110;
DRAM[61304] = 8'b1111101;
DRAM[61305] = 8'b10000010;
DRAM[61306] = 8'b1101110;
DRAM[61307] = 8'b1110000;
DRAM[61308] = 8'b1111011;
DRAM[61309] = 8'b1110111;
DRAM[61310] = 8'b1110101;
DRAM[61311] = 8'b1101100;
DRAM[61312] = 8'b1101011;
DRAM[61313] = 8'b1100111;
DRAM[61314] = 8'b1101111;
DRAM[61315] = 8'b1101001;
DRAM[61316] = 8'b1101101;
DRAM[61317] = 8'b1111001;
DRAM[61318] = 8'b1101111;
DRAM[61319] = 8'b1110000;
DRAM[61320] = 8'b1111000;
DRAM[61321] = 8'b1101101;
DRAM[61322] = 8'b1101100;
DRAM[61323] = 8'b1110110;
DRAM[61324] = 8'b1110100;
DRAM[61325] = 8'b1101001;
DRAM[61326] = 8'b1101011;
DRAM[61327] = 8'b1110111;
DRAM[61328] = 8'b1101000;
DRAM[61329] = 8'b1111000;
DRAM[61330] = 8'b1101101;
DRAM[61331] = 8'b1100101;
DRAM[61332] = 8'b1110101;
DRAM[61333] = 8'b1101101;
DRAM[61334] = 8'b1100001;
DRAM[61335] = 8'b1110001;
DRAM[61336] = 8'b1111001;
DRAM[61337] = 8'b1110011;
DRAM[61338] = 8'b1101111;
DRAM[61339] = 8'b1110010;
DRAM[61340] = 8'b1110110;
DRAM[61341] = 8'b1111000;
DRAM[61342] = 8'b1110110;
DRAM[61343] = 8'b1110101;
DRAM[61344] = 8'b10001101;
DRAM[61345] = 8'b1111011;
DRAM[61346] = 8'b1110110;
DRAM[61347] = 8'b1101010;
DRAM[61348] = 8'b1110000;
DRAM[61349] = 8'b10000000;
DRAM[61350] = 8'b10000001;
DRAM[61351] = 8'b10001011;
DRAM[61352] = 8'b10000111;
DRAM[61353] = 8'b10001101;
DRAM[61354] = 8'b10010011;
DRAM[61355] = 8'b10010101;
DRAM[61356] = 8'b10010101;
DRAM[61357] = 8'b10011000;
DRAM[61358] = 8'b10100001;
DRAM[61359] = 8'b10101000;
DRAM[61360] = 8'b10011011;
DRAM[61361] = 8'b10011100;
DRAM[61362] = 8'b10100010;
DRAM[61363] = 8'b10101011;
DRAM[61364] = 8'b10110000;
DRAM[61365] = 8'b10110010;
DRAM[61366] = 8'b10110111;
DRAM[61367] = 8'b10111101;
DRAM[61368] = 8'b10111110;
DRAM[61369] = 8'b11000011;
DRAM[61370] = 8'b11001100;
DRAM[61371] = 8'b11011001;
DRAM[61372] = 8'b11100101;
DRAM[61373] = 8'b11101100;
DRAM[61374] = 8'b11101111;
DRAM[61375] = 8'b11101111;
DRAM[61376] = 8'b11110111;
DRAM[61377] = 8'b11101001;
DRAM[61378] = 8'b11010101;
DRAM[61379] = 8'b11000001;
DRAM[61380] = 8'b10101111;
DRAM[61381] = 8'b10100000;
DRAM[61382] = 8'b10011000;
DRAM[61383] = 8'b10010110;
DRAM[61384] = 8'b10011001;
DRAM[61385] = 8'b10011000;
DRAM[61386] = 8'b10010101;
DRAM[61387] = 8'b10010001;
DRAM[61388] = 8'b10001100;
DRAM[61389] = 8'b10001000;
DRAM[61390] = 8'b10000100;
DRAM[61391] = 8'b10000001;
DRAM[61392] = 8'b1111011;
DRAM[61393] = 8'b1111010;
DRAM[61394] = 8'b1111001;
DRAM[61395] = 8'b1110111;
DRAM[61396] = 8'b1110101;
DRAM[61397] = 8'b1110011;
DRAM[61398] = 8'b1110010;
DRAM[61399] = 8'b1110001;
DRAM[61400] = 8'b1101111;
DRAM[61401] = 8'b1101111;
DRAM[61402] = 8'b1101111;
DRAM[61403] = 8'b1101110;
DRAM[61404] = 8'b1101101;
DRAM[61405] = 8'b1101101;
DRAM[61406] = 8'b1101100;
DRAM[61407] = 8'b1101100;
DRAM[61408] = 8'b1101010;
DRAM[61409] = 8'b1101001;
DRAM[61410] = 8'b1101000;
DRAM[61411] = 8'b1100111;
DRAM[61412] = 8'b1100111;
DRAM[61413] = 8'b1100111;
DRAM[61414] = 8'b1100111;
DRAM[61415] = 8'b1101000;
DRAM[61416] = 8'b1101000;
DRAM[61417] = 8'b1100111;
DRAM[61418] = 8'b1100111;
DRAM[61419] = 8'b1100111;
DRAM[61420] = 8'b1100111;
DRAM[61421] = 8'b1101000;
DRAM[61422] = 8'b1101001;
DRAM[61423] = 8'b1101010;
DRAM[61424] = 8'b1101010;
DRAM[61425] = 8'b1101011;
DRAM[61426] = 8'b1101101;
DRAM[61427] = 8'b1110000;
DRAM[61428] = 8'b1110010;
DRAM[61429] = 8'b1110010;
DRAM[61430] = 8'b1101111;
DRAM[61431] = 8'b1101100;
DRAM[61432] = 8'b1101100;
DRAM[61433] = 8'b1101100;
DRAM[61434] = 8'b1101100;
DRAM[61435] = 8'b1101011;
DRAM[61436] = 8'b1101010;
DRAM[61437] = 8'b1101001;
DRAM[61438] = 8'b1100111;
DRAM[61439] = 8'b1100110;
DRAM[61440] = 8'b10010001;
DRAM[61441] = 8'b10010001;
DRAM[61442] = 8'b10010000;
DRAM[61443] = 8'b10001110;
DRAM[61444] = 8'b10001110;
DRAM[61445] = 8'b10001110;
DRAM[61446] = 8'b10001100;
DRAM[61447] = 8'b10001000;
DRAM[61448] = 8'b10010011;
DRAM[61449] = 8'b10011010;
DRAM[61450] = 8'b10101010;
DRAM[61451] = 8'b11000011;
DRAM[61452] = 8'b11100001;
DRAM[61453] = 8'b11110110;
DRAM[61454] = 8'b11111000;
DRAM[61455] = 8'b11110000;
DRAM[61456] = 8'b11111001;
DRAM[61457] = 8'b11110110;
DRAM[61458] = 8'b11110010;
DRAM[61459] = 8'b11110010;
DRAM[61460] = 8'b11110100;
DRAM[61461] = 8'b11110100;
DRAM[61462] = 8'b11110001;
DRAM[61463] = 8'b11101101;
DRAM[61464] = 8'b11110001;
DRAM[61465] = 8'b11101111;
DRAM[61466] = 8'b11101101;
DRAM[61467] = 8'b11101001;
DRAM[61468] = 8'b11100110;
DRAM[61469] = 8'b11100011;
DRAM[61470] = 8'b11100000;
DRAM[61471] = 8'b11011111;
DRAM[61472] = 8'b11011010;
DRAM[61473] = 8'b11010001;
DRAM[61474] = 8'b11001000;
DRAM[61475] = 8'b11000111;
DRAM[61476] = 8'b11001100;
DRAM[61477] = 8'b11001101;
DRAM[61478] = 8'b11001001;
DRAM[61479] = 8'b11000011;
DRAM[61480] = 8'b11001000;
DRAM[61481] = 8'b10111110;
DRAM[61482] = 8'b10110100;
DRAM[61483] = 8'b10110011;
DRAM[61484] = 8'b10110101;
DRAM[61485] = 8'b10110011;
DRAM[61486] = 8'b10101000;
DRAM[61487] = 8'b10011101;
DRAM[61488] = 8'b10101001;
DRAM[61489] = 8'b10100100;
DRAM[61490] = 8'b10011111;
DRAM[61491] = 8'b10011110;
DRAM[61492] = 8'b10100001;
DRAM[61493] = 8'b10100011;
DRAM[61494] = 8'b10100010;
DRAM[61495] = 8'b10100000;
DRAM[61496] = 8'b10011111;
DRAM[61497] = 8'b10101001;
DRAM[61498] = 8'b10101101;
DRAM[61499] = 8'b10100110;
DRAM[61500] = 8'b10011111;
DRAM[61501] = 8'b10011100;
DRAM[61502] = 8'b10011010;
DRAM[61503] = 8'b10010110;
DRAM[61504] = 8'b10000110;
DRAM[61505] = 8'b1111101;
DRAM[61506] = 8'b1111000;
DRAM[61507] = 8'b1110110;
DRAM[61508] = 8'b1110000;
DRAM[61509] = 8'b1101100;
DRAM[61510] = 8'b1110111;
DRAM[61511] = 8'b10000111;
DRAM[61512] = 8'b10001101;
DRAM[61513] = 8'b10011001;
DRAM[61514] = 8'b10011011;
DRAM[61515] = 8'b10001101;
DRAM[61516] = 8'b10000010;
DRAM[61517] = 8'b10000011;
DRAM[61518] = 8'b10000011;
DRAM[61519] = 8'b1111110;
DRAM[61520] = 8'b1111010;
DRAM[61521] = 8'b1111100;
DRAM[61522] = 8'b10001111;
DRAM[61523] = 8'b1111100;
DRAM[61524] = 8'b1110101;
DRAM[61525] = 8'b10000011;
DRAM[61526] = 8'b1110110;
DRAM[61527] = 8'b1111111;
DRAM[61528] = 8'b1101110;
DRAM[61529] = 8'b10000101;
DRAM[61530] = 8'b10001101;
DRAM[61531] = 8'b1111100;
DRAM[61532] = 8'b1110010;
DRAM[61533] = 8'b1111010;
DRAM[61534] = 8'b1111101;
DRAM[61535] = 8'b1110101;
DRAM[61536] = 8'b1110100;
DRAM[61537] = 8'b1101000;
DRAM[61538] = 8'b1101111;
DRAM[61539] = 8'b1111100;
DRAM[61540] = 8'b1110110;
DRAM[61541] = 8'b1101100;
DRAM[61542] = 8'b1101100;
DRAM[61543] = 8'b1101011;
DRAM[61544] = 8'b1110010;
DRAM[61545] = 8'b1111010;
DRAM[61546] = 8'b1111100;
DRAM[61547] = 8'b1110000;
DRAM[61548] = 8'b1100010;
DRAM[61549] = 8'b1100000;
DRAM[61550] = 8'b1101010;
DRAM[61551] = 8'b1110101;
DRAM[61552] = 8'b1101010;
DRAM[61553] = 8'b1100111;
DRAM[61554] = 8'b1101101;
DRAM[61555] = 8'b1110100;
DRAM[61556] = 8'b1101110;
DRAM[61557] = 8'b1100010;
DRAM[61558] = 8'b1101001;
DRAM[61559] = 8'b1111010;
DRAM[61560] = 8'b1111001;
DRAM[61561] = 8'b10000001;
DRAM[61562] = 8'b1110001;
DRAM[61563] = 8'b1101011;
DRAM[61564] = 8'b1101011;
DRAM[61565] = 8'b1110000;
DRAM[61566] = 8'b1111101;
DRAM[61567] = 8'b1110011;
DRAM[61568] = 8'b1100011;
DRAM[61569] = 8'b1101110;
DRAM[61570] = 8'b1110100;
DRAM[61571] = 8'b1110000;
DRAM[61572] = 8'b1101011;
DRAM[61573] = 8'b1101101;
DRAM[61574] = 8'b1101110;
DRAM[61575] = 8'b1101100;
DRAM[61576] = 8'b1101100;
DRAM[61577] = 8'b1101110;
DRAM[61578] = 8'b1110001;
DRAM[61579] = 8'b1110000;
DRAM[61580] = 8'b1101010;
DRAM[61581] = 8'b1100110;
DRAM[61582] = 8'b1101001;
DRAM[61583] = 8'b1101110;
DRAM[61584] = 8'b1110000;
DRAM[61585] = 8'b1110110;
DRAM[61586] = 8'b1101101;
DRAM[61587] = 8'b1100100;
DRAM[61588] = 8'b1101100;
DRAM[61589] = 8'b1110010;
DRAM[61590] = 8'b1110000;
DRAM[61591] = 8'b1110000;
DRAM[61592] = 8'b1110010;
DRAM[61593] = 8'b1110010;
DRAM[61594] = 8'b1110000;
DRAM[61595] = 8'b1101111;
DRAM[61596] = 8'b1110010;
DRAM[61597] = 8'b1110111;
DRAM[61598] = 8'b1110101;
DRAM[61599] = 8'b1110000;
DRAM[61600] = 8'b1111011;
DRAM[61601] = 8'b1111111;
DRAM[61602] = 8'b10000010;
DRAM[61603] = 8'b1111110;
DRAM[61604] = 8'b1111001;
DRAM[61605] = 8'b1111000;
DRAM[61606] = 8'b1111111;
DRAM[61607] = 8'b10000110;
DRAM[61608] = 8'b10000101;
DRAM[61609] = 8'b10001101;
DRAM[61610] = 8'b10001111;
DRAM[61611] = 8'b10001100;
DRAM[61612] = 8'b10010001;
DRAM[61613] = 8'b10011110;
DRAM[61614] = 8'b10100100;
DRAM[61615] = 8'b10100010;
DRAM[61616] = 8'b10100001;
DRAM[61617] = 8'b10100101;
DRAM[61618] = 8'b10101100;
DRAM[61619] = 8'b10110010;
DRAM[61620] = 8'b10110101;
DRAM[61621] = 8'b10110110;
DRAM[61622] = 8'b10110101;
DRAM[61623] = 8'b10110100;
DRAM[61624] = 8'b11000000;
DRAM[61625] = 8'b11000111;
DRAM[61626] = 8'b11001011;
DRAM[61627] = 8'b11001011;
DRAM[61628] = 8'b11010010;
DRAM[61629] = 8'b11100001;
DRAM[61630] = 8'b11101011;
DRAM[61631] = 8'b11101110;
DRAM[61632] = 8'b11110100;
DRAM[61633] = 8'b11111000;
DRAM[61634] = 8'b11101101;
DRAM[61635] = 8'b11010010;
DRAM[61636] = 8'b10111010;
DRAM[61637] = 8'b10101101;
DRAM[61638] = 8'b10100110;
DRAM[61639] = 8'b10100000;
DRAM[61640] = 8'b10011100;
DRAM[61641] = 8'b10011001;
DRAM[61642] = 8'b10010110;
DRAM[61643] = 8'b10010011;
DRAM[61644] = 8'b10010010;
DRAM[61645] = 8'b10001111;
DRAM[61646] = 8'b10001100;
DRAM[61647] = 8'b10001001;
DRAM[61648] = 8'b1111010;
DRAM[61649] = 8'b1111001;
DRAM[61650] = 8'b1111000;
DRAM[61651] = 8'b1110101;
DRAM[61652] = 8'b1110010;
DRAM[61653] = 8'b1101111;
DRAM[61654] = 8'b1101101;
DRAM[61655] = 8'b1101011;
DRAM[61656] = 8'b1101111;
DRAM[61657] = 8'b1101111;
DRAM[61658] = 8'b1101110;
DRAM[61659] = 8'b1101110;
DRAM[61660] = 8'b1101101;
DRAM[61661] = 8'b1101100;
DRAM[61662] = 8'b1101100;
DRAM[61663] = 8'b1101011;
DRAM[61664] = 8'b1100111;
DRAM[61665] = 8'b1100111;
DRAM[61666] = 8'b1100111;
DRAM[61667] = 8'b1100111;
DRAM[61668] = 8'b1100111;
DRAM[61669] = 8'b1100111;
DRAM[61670] = 8'b1100111;
DRAM[61671] = 8'b1100111;
DRAM[61672] = 8'b1101001;
DRAM[61673] = 8'b1101000;
DRAM[61674] = 8'b1101000;
DRAM[61675] = 8'b1100111;
DRAM[61676] = 8'b1100111;
DRAM[61677] = 8'b1101000;
DRAM[61678] = 8'b1101000;
DRAM[61679] = 8'b1101001;
DRAM[61680] = 8'b1101011;
DRAM[61681] = 8'b1101100;
DRAM[61682] = 8'b1101111;
DRAM[61683] = 8'b1110001;
DRAM[61684] = 8'b1110010;
DRAM[61685] = 8'b1110001;
DRAM[61686] = 8'b1110000;
DRAM[61687] = 8'b1101111;
DRAM[61688] = 8'b1101100;
DRAM[61689] = 8'b1101100;
DRAM[61690] = 8'b1101011;
DRAM[61691] = 8'b1101010;
DRAM[61692] = 8'b1101001;
DRAM[61693] = 8'b1100111;
DRAM[61694] = 8'b1100111;
DRAM[61695] = 8'b1100110;
DRAM[61696] = 8'b10010001;
DRAM[61697] = 8'b10010000;
DRAM[61698] = 8'b10001111;
DRAM[61699] = 8'b10001101;
DRAM[61700] = 8'b10001101;
DRAM[61701] = 8'b10001100;
DRAM[61702] = 8'b10001011;
DRAM[61703] = 8'b10001001;
DRAM[61704] = 8'b10010101;
DRAM[61705] = 8'b10100110;
DRAM[61706] = 8'b10111101;
DRAM[61707] = 8'b11010101;
DRAM[61708] = 8'b11101011;
DRAM[61709] = 8'b11111010;
DRAM[61710] = 8'b11111100;
DRAM[61711] = 8'b11110111;
DRAM[61712] = 8'b11110111;
DRAM[61713] = 8'b11110100;
DRAM[61714] = 8'b11110010;
DRAM[61715] = 8'b11110010;
DRAM[61716] = 8'b11110100;
DRAM[61717] = 8'b11110100;
DRAM[61718] = 8'b11110001;
DRAM[61719] = 8'b11101101;
DRAM[61720] = 8'b11101001;
DRAM[61721] = 8'b11100110;
DRAM[61722] = 8'b11100011;
DRAM[61723] = 8'b11100010;
DRAM[61724] = 8'b11100001;
DRAM[61725] = 8'b11100000;
DRAM[61726] = 8'b11011101;
DRAM[61727] = 8'b11011010;
DRAM[61728] = 8'b11010000;
DRAM[61729] = 8'b11001001;
DRAM[61730] = 8'b11000010;
DRAM[61731] = 8'b11000011;
DRAM[61732] = 8'b11000111;
DRAM[61733] = 8'b11001010;
DRAM[61734] = 8'b11000110;
DRAM[61735] = 8'b11000000;
DRAM[61736] = 8'b10111011;
DRAM[61737] = 8'b10111010;
DRAM[61738] = 8'b10110111;
DRAM[61739] = 8'b10110000;
DRAM[61740] = 8'b10101010;
DRAM[61741] = 8'b10100110;
DRAM[61742] = 8'b10100111;
DRAM[61743] = 8'b10101001;
DRAM[61744] = 8'b10100111;
DRAM[61745] = 8'b10100111;
DRAM[61746] = 8'b10100101;
DRAM[61747] = 8'b10100000;
DRAM[61748] = 8'b10011010;
DRAM[61749] = 8'b10010101;
DRAM[61750] = 8'b10010001;
DRAM[61751] = 8'b10001111;
DRAM[61752] = 8'b10010101;
DRAM[61753] = 8'b10011010;
DRAM[61754] = 8'b10011011;
DRAM[61755] = 8'b10010100;
DRAM[61756] = 8'b10001110;
DRAM[61757] = 8'b10001110;
DRAM[61758] = 8'b10001101;
DRAM[61759] = 8'b10001011;
DRAM[61760] = 8'b10001100;
DRAM[61761] = 8'b10000110;
DRAM[61762] = 8'b10000000;
DRAM[61763] = 8'b1111000;
DRAM[61764] = 8'b1101111;
DRAM[61765] = 8'b1101001;
DRAM[61766] = 8'b1101011;
DRAM[61767] = 8'b1110001;
DRAM[61768] = 8'b10000000;
DRAM[61769] = 8'b10000101;
DRAM[61770] = 8'b10001100;
DRAM[61771] = 8'b10001110;
DRAM[61772] = 8'b10001001;
DRAM[61773] = 8'b10000100;
DRAM[61774] = 8'b10000110;
DRAM[61775] = 8'b10001011;
DRAM[61776] = 8'b10000011;
DRAM[61777] = 8'b10000101;
DRAM[61778] = 8'b10001101;
DRAM[61779] = 8'b10000100;
DRAM[61780] = 8'b1111101;
DRAM[61781] = 8'b1111110;
DRAM[61782] = 8'b1110110;
DRAM[61783] = 8'b1111000;
DRAM[61784] = 8'b1111110;
DRAM[61785] = 8'b1111000;
DRAM[61786] = 8'b1110100;
DRAM[61787] = 8'b1111000;
DRAM[61788] = 8'b10000000;
DRAM[61789] = 8'b10000100;
DRAM[61790] = 8'b1111101;
DRAM[61791] = 8'b1110011;
DRAM[61792] = 8'b1110010;
DRAM[61793] = 8'b1110110;
DRAM[61794] = 8'b1111100;
DRAM[61795] = 8'b1110100;
DRAM[61796] = 8'b1101011;
DRAM[61797] = 8'b1110001;
DRAM[61798] = 8'b1110011;
DRAM[61799] = 8'b1100100;
DRAM[61800] = 8'b1110010;
DRAM[61801] = 8'b1100110;
DRAM[61802] = 8'b1101100;
DRAM[61803] = 8'b10000000;
DRAM[61804] = 8'b1111110;
DRAM[61805] = 8'b1100110;
DRAM[61806] = 8'b1011101;
DRAM[61807] = 8'b1101000;
DRAM[61808] = 8'b1110001;
DRAM[61809] = 8'b1100000;
DRAM[61810] = 8'b1011000;
DRAM[61811] = 8'b1100101;
DRAM[61812] = 8'b1110100;
DRAM[61813] = 8'b1110010;
DRAM[61814] = 8'b1100110;
DRAM[61815] = 8'b1011110;
DRAM[61816] = 8'b1101000;
DRAM[61817] = 8'b1110101;
DRAM[61818] = 8'b1110011;
DRAM[61819] = 8'b1111001;
DRAM[61820] = 8'b1110010;
DRAM[61821] = 8'b1100111;
DRAM[61822] = 8'b1110110;
DRAM[61823] = 8'b1111001;
DRAM[61824] = 8'b1011100;
DRAM[61825] = 8'b1101001;
DRAM[61826] = 8'b1110010;
DRAM[61827] = 8'b1101111;
DRAM[61828] = 8'b1101011;
DRAM[61829] = 8'b1110000;
DRAM[61830] = 8'b1111000;
DRAM[61831] = 8'b1111100;
DRAM[61832] = 8'b1101001;
DRAM[61833] = 8'b1101010;
DRAM[61834] = 8'b1101100;
DRAM[61835] = 8'b1101100;
DRAM[61836] = 8'b1101010;
DRAM[61837] = 8'b1101001;
DRAM[61838] = 8'b1101011;
DRAM[61839] = 8'b1101110;
DRAM[61840] = 8'b1101001;
DRAM[61841] = 8'b1110000;
DRAM[61842] = 8'b1101010;
DRAM[61843] = 8'b1100011;
DRAM[61844] = 8'b1100111;
DRAM[61845] = 8'b1101000;
DRAM[61846] = 8'b1101000;
DRAM[61847] = 8'b1101111;
DRAM[61848] = 8'b1110001;
DRAM[61849] = 8'b1110011;
DRAM[61850] = 8'b1110010;
DRAM[61851] = 8'b1101101;
DRAM[61852] = 8'b1101101;
DRAM[61853] = 8'b1110010;
DRAM[61854] = 8'b1110111;
DRAM[61855] = 8'b1111000;
DRAM[61856] = 8'b1111010;
DRAM[61857] = 8'b1111111;
DRAM[61858] = 8'b10000010;
DRAM[61859] = 8'b1111111;
DRAM[61860] = 8'b1111010;
DRAM[61861] = 8'b1111001;
DRAM[61862] = 8'b1111111;
DRAM[61863] = 8'b10000100;
DRAM[61864] = 8'b10000100;
DRAM[61865] = 8'b10001101;
DRAM[61866] = 8'b10010101;
DRAM[61867] = 8'b10010101;
DRAM[61868] = 8'b10010100;
DRAM[61869] = 8'b10011000;
DRAM[61870] = 8'b10011101;
DRAM[61871] = 8'b10100000;
DRAM[61872] = 8'b10011100;
DRAM[61873] = 8'b10011110;
DRAM[61874] = 8'b10100010;
DRAM[61875] = 8'b10101001;
DRAM[61876] = 8'b10110010;
DRAM[61877] = 8'b10111000;
DRAM[61878] = 8'b10111010;
DRAM[61879] = 8'b10111001;
DRAM[61880] = 8'b10111001;
DRAM[61881] = 8'b11000000;
DRAM[61882] = 8'b11000110;
DRAM[61883] = 8'b11001001;
DRAM[61884] = 8'b11010001;
DRAM[61885] = 8'b11100000;
DRAM[61886] = 8'b11101011;
DRAM[61887] = 8'b11101110;
DRAM[61888] = 8'b11110010;
DRAM[61889] = 8'b11110101;
DRAM[61890] = 8'b11101100;
DRAM[61891] = 8'b11011000;
DRAM[61892] = 8'b11000111;
DRAM[61893] = 8'b10111101;
DRAM[61894] = 8'b10110001;
DRAM[61895] = 8'b10100101;
DRAM[61896] = 8'b10011101;
DRAM[61897] = 8'b10011010;
DRAM[61898] = 8'b10010101;
DRAM[61899] = 8'b10010001;
DRAM[61900] = 8'b10001101;
DRAM[61901] = 8'b10001001;
DRAM[61902] = 8'b10000101;
DRAM[61903] = 8'b10000001;
DRAM[61904] = 8'b1111001;
DRAM[61905] = 8'b1111001;
DRAM[61906] = 8'b1110111;
DRAM[61907] = 8'b1110101;
DRAM[61908] = 8'b1110010;
DRAM[61909] = 8'b1101111;
DRAM[61910] = 8'b1101100;
DRAM[61911] = 8'b1101011;
DRAM[61912] = 8'b1101110;
DRAM[61913] = 8'b1101101;
DRAM[61914] = 8'b1101101;
DRAM[61915] = 8'b1101101;
DRAM[61916] = 8'b1101100;
DRAM[61917] = 8'b1101011;
DRAM[61918] = 8'b1101011;
DRAM[61919] = 8'b1101011;
DRAM[61920] = 8'b1100111;
DRAM[61921] = 8'b1100111;
DRAM[61922] = 8'b1100111;
DRAM[61923] = 8'b1100111;
DRAM[61924] = 8'b1100111;
DRAM[61925] = 8'b1100111;
DRAM[61926] = 8'b1100111;
DRAM[61927] = 8'b1100111;
DRAM[61928] = 8'b1101001;
DRAM[61929] = 8'b1101000;
DRAM[61930] = 8'b1101000;
DRAM[61931] = 8'b1100111;
DRAM[61932] = 8'b1100111;
DRAM[61933] = 8'b1101000;
DRAM[61934] = 8'b1101000;
DRAM[61935] = 8'b1101001;
DRAM[61936] = 8'b1101010;
DRAM[61937] = 8'b1101100;
DRAM[61938] = 8'b1101111;
DRAM[61939] = 8'b1110001;
DRAM[61940] = 8'b1110010;
DRAM[61941] = 8'b1110001;
DRAM[61942] = 8'b1110000;
DRAM[61943] = 8'b1101111;
DRAM[61944] = 8'b1101100;
DRAM[61945] = 8'b1101011;
DRAM[61946] = 8'b1101010;
DRAM[61947] = 8'b1101001;
DRAM[61948] = 8'b1101000;
DRAM[61949] = 8'b1100111;
DRAM[61950] = 8'b1100110;
DRAM[61951] = 8'b1100101;
DRAM[61952] = 8'b10010000;
DRAM[61953] = 8'b10001111;
DRAM[61954] = 8'b10001101;
DRAM[61955] = 8'b10001100;
DRAM[61956] = 8'b10001011;
DRAM[61957] = 8'b10001010;
DRAM[61958] = 8'b10001010;
DRAM[61959] = 8'b10001011;
DRAM[61960] = 8'b10010011;
DRAM[61961] = 8'b10101101;
DRAM[61962] = 8'b11001100;
DRAM[61963] = 8'b11100010;
DRAM[61964] = 8'b11101110;
DRAM[61965] = 8'b11110101;
DRAM[61966] = 8'b11110111;
DRAM[61967] = 8'b11110101;
DRAM[61968] = 8'b11110101;
DRAM[61969] = 8'b11110010;
DRAM[61970] = 8'b11110000;
DRAM[61971] = 8'b11110001;
DRAM[61972] = 8'b11110100;
DRAM[61973] = 8'b11110100;
DRAM[61974] = 8'b11110001;
DRAM[61975] = 8'b11101101;
DRAM[61976] = 8'b11100111;
DRAM[61977] = 8'b11100011;
DRAM[61978] = 8'b11011110;
DRAM[61979] = 8'b11011111;
DRAM[61980] = 8'b11100010;
DRAM[61981] = 8'b11100010;
DRAM[61982] = 8'b11011110;
DRAM[61983] = 8'b11011001;
DRAM[61984] = 8'b11010101;
DRAM[61985] = 8'b11010000;
DRAM[61986] = 8'b11001101;
DRAM[61987] = 8'b11001110;
DRAM[61988] = 8'b11010011;
DRAM[61989] = 8'b11010100;
DRAM[61990] = 8'b11010001;
DRAM[61991] = 8'b11001101;
DRAM[61992] = 8'b11000111;
DRAM[61993] = 8'b11000101;
DRAM[61994] = 8'b11000000;
DRAM[61995] = 8'b10111001;
DRAM[61996] = 8'b10110011;
DRAM[61997] = 8'b10110010;
DRAM[61998] = 8'b10110101;
DRAM[61999] = 8'b10111001;
DRAM[62000] = 8'b10101011;
DRAM[62001] = 8'b10101100;
DRAM[62002] = 8'b10101011;
DRAM[62003] = 8'b10100100;
DRAM[62004] = 8'b10011011;
DRAM[62005] = 8'b10010110;
DRAM[62006] = 8'b10010110;
DRAM[62007] = 8'b10011001;
DRAM[62008] = 8'b10010100;
DRAM[62009] = 8'b10011000;
DRAM[62010] = 8'b10011001;
DRAM[62011] = 8'b10010111;
DRAM[62012] = 8'b10010101;
DRAM[62013] = 8'b10010100;
DRAM[62014] = 8'b10010001;
DRAM[62015] = 8'b10001101;
DRAM[62016] = 8'b10001100;
DRAM[62017] = 8'b10001101;
DRAM[62018] = 8'b10001001;
DRAM[62019] = 8'b10000001;
DRAM[62020] = 8'b1111100;
DRAM[62021] = 8'b1111010;
DRAM[62022] = 8'b1110111;
DRAM[62023] = 8'b1110011;
DRAM[62024] = 8'b1111001;
DRAM[62025] = 8'b1110110;
DRAM[62026] = 8'b1111111;
DRAM[62027] = 8'b10001110;
DRAM[62028] = 8'b10010010;
DRAM[62029] = 8'b10001010;
DRAM[62030] = 8'b10001100;
DRAM[62031] = 8'b10010110;
DRAM[62032] = 8'b10000100;
DRAM[62033] = 8'b10000111;
DRAM[62034] = 8'b10000010;
DRAM[62035] = 8'b10001001;
DRAM[62036] = 8'b10001000;
DRAM[62037] = 8'b1111110;
DRAM[62038] = 8'b10000001;
DRAM[62039] = 8'b1111101;
DRAM[62040] = 8'b10001001;
DRAM[62041] = 8'b1110001;
DRAM[62042] = 8'b1101000;
DRAM[62043] = 8'b1111010;
DRAM[62044] = 8'b10001000;
DRAM[62045] = 8'b10000010;
DRAM[62046] = 8'b1110111;
DRAM[62047] = 8'b1110110;
DRAM[62048] = 8'b1110010;
DRAM[62049] = 8'b1110111;
DRAM[62050] = 8'b1111100;
DRAM[62051] = 8'b1110100;
DRAM[62052] = 8'b1101100;
DRAM[62053] = 8'b1110011;
DRAM[62054] = 8'b1110110;
DRAM[62055] = 8'b1100111;
DRAM[62056] = 8'b1101100;
DRAM[62057] = 8'b1110011;
DRAM[62058] = 8'b1110101;
DRAM[62059] = 8'b1110001;
DRAM[62060] = 8'b1101111;
DRAM[62061] = 8'b1110000;
DRAM[62062] = 8'b1101001;
DRAM[62063] = 8'b1011111;
DRAM[62064] = 8'b1101100;
DRAM[62065] = 8'b1100011;
DRAM[62066] = 8'b1011100;
DRAM[62067] = 8'b1100001;
DRAM[62068] = 8'b1101101;
DRAM[62069] = 8'b1110100;
DRAM[62070] = 8'b1110001;
DRAM[62071] = 8'b1101011;
DRAM[62072] = 8'b1100001;
DRAM[62073] = 8'b1101000;
DRAM[62074] = 8'b1101011;
DRAM[62075] = 8'b1111101;
DRAM[62076] = 8'b1111001;
DRAM[62077] = 8'b1100110;
DRAM[62078] = 8'b1101110;
DRAM[62079] = 8'b1110100;
DRAM[62080] = 8'b1100100;
DRAM[62081] = 8'b1101111;
DRAM[62082] = 8'b1110110;
DRAM[62083] = 8'b1110001;
DRAM[62084] = 8'b1101010;
DRAM[62085] = 8'b1101100;
DRAM[62086] = 8'b1110100;
DRAM[62087] = 8'b1111011;
DRAM[62088] = 8'b1101000;
DRAM[62089] = 8'b1101000;
DRAM[62090] = 8'b1100111;
DRAM[62091] = 8'b1100111;
DRAM[62092] = 8'b1101001;
DRAM[62093] = 8'b1101011;
DRAM[62094] = 8'b1101100;
DRAM[62095] = 8'b1101011;
DRAM[62096] = 8'b1100110;
DRAM[62097] = 8'b1101011;
DRAM[62098] = 8'b1101000;
DRAM[62099] = 8'b1100101;
DRAM[62100] = 8'b1100111;
DRAM[62101] = 8'b1100010;
DRAM[62102] = 8'b1100011;
DRAM[62103] = 8'b1110000;
DRAM[62104] = 8'b1101101;
DRAM[62105] = 8'b1110010;
DRAM[62106] = 8'b1110001;
DRAM[62107] = 8'b1101010;
DRAM[62108] = 8'b1100110;
DRAM[62109] = 8'b1101100;
DRAM[62110] = 8'b1110110;
DRAM[62111] = 8'b1111101;
DRAM[62112] = 8'b1111001;
DRAM[62113] = 8'b1111110;
DRAM[62114] = 8'b10000010;
DRAM[62115] = 8'b10000001;
DRAM[62116] = 8'b1111101;
DRAM[62117] = 8'b1111011;
DRAM[62118] = 8'b1111110;
DRAM[62119] = 8'b10000010;
DRAM[62120] = 8'b10000011;
DRAM[62121] = 8'b10001011;
DRAM[62122] = 8'b10010111;
DRAM[62123] = 8'b10011100;
DRAM[62124] = 8'b10011000;
DRAM[62125] = 8'b10010010;
DRAM[62126] = 8'b10010110;
DRAM[62127] = 8'b10011101;
DRAM[62128] = 8'b10100011;
DRAM[62129] = 8'b10100010;
DRAM[62130] = 8'b10100100;
DRAM[62131] = 8'b10101010;
DRAM[62132] = 8'b10110011;
DRAM[62133] = 8'b10111011;
DRAM[62134] = 8'b10111111;
DRAM[62135] = 8'b10111111;
DRAM[62136] = 8'b10111111;
DRAM[62137] = 8'b11000100;
DRAM[62138] = 8'b11000111;
DRAM[62139] = 8'b11001001;
DRAM[62140] = 8'b11001101;
DRAM[62141] = 8'b11010111;
DRAM[62142] = 8'b11011110;
DRAM[62143] = 8'b11100001;
DRAM[62144] = 8'b11110011;
DRAM[62145] = 8'b11110000;
DRAM[62146] = 8'b11100100;
DRAM[62147] = 8'b11010000;
DRAM[62148] = 8'b11000011;
DRAM[62149] = 8'b10111011;
DRAM[62150] = 8'b10101101;
DRAM[62151] = 8'b10011110;
DRAM[62152] = 8'b10011001;
DRAM[62153] = 8'b10010110;
DRAM[62154] = 8'b10010001;
DRAM[62155] = 8'b10001100;
DRAM[62156] = 8'b10001000;
DRAM[62157] = 8'b10000100;
DRAM[62158] = 8'b1111111;
DRAM[62159] = 8'b1111011;
DRAM[62160] = 8'b1111000;
DRAM[62161] = 8'b1110111;
DRAM[62162] = 8'b1110110;
DRAM[62163] = 8'b1110100;
DRAM[62164] = 8'b1110001;
DRAM[62165] = 8'b1101110;
DRAM[62166] = 8'b1101011;
DRAM[62167] = 8'b1101001;
DRAM[62168] = 8'b1101011;
DRAM[62169] = 8'b1101011;
DRAM[62170] = 8'b1101011;
DRAM[62171] = 8'b1101011;
DRAM[62172] = 8'b1101010;
DRAM[62173] = 8'b1101010;
DRAM[62174] = 8'b1101010;
DRAM[62175] = 8'b1101010;
DRAM[62176] = 8'b1100110;
DRAM[62177] = 8'b1100110;
DRAM[62178] = 8'b1100110;
DRAM[62179] = 8'b1100111;
DRAM[62180] = 8'b1100111;
DRAM[62181] = 8'b1100111;
DRAM[62182] = 8'b1100111;
DRAM[62183] = 8'b1100111;
DRAM[62184] = 8'b1101001;
DRAM[62185] = 8'b1101000;
DRAM[62186] = 8'b1101000;
DRAM[62187] = 8'b1100111;
DRAM[62188] = 8'b1100111;
DRAM[62189] = 8'b1101000;
DRAM[62190] = 8'b1101000;
DRAM[62191] = 8'b1101001;
DRAM[62192] = 8'b1101010;
DRAM[62193] = 8'b1101100;
DRAM[62194] = 8'b1101110;
DRAM[62195] = 8'b1110001;
DRAM[62196] = 8'b1110001;
DRAM[62197] = 8'b1110001;
DRAM[62198] = 8'b1101111;
DRAM[62199] = 8'b1101110;
DRAM[62200] = 8'b1101011;
DRAM[62201] = 8'b1101010;
DRAM[62202] = 8'b1101001;
DRAM[62203] = 8'b1101000;
DRAM[62204] = 8'b1100111;
DRAM[62205] = 8'b1100110;
DRAM[62206] = 8'b1100101;
DRAM[62207] = 8'b1100100;
DRAM[62208] = 8'b10010000;
DRAM[62209] = 8'b10001101;
DRAM[62210] = 8'b10001011;
DRAM[62211] = 8'b10001011;
DRAM[62212] = 8'b10001001;
DRAM[62213] = 8'b10001000;
DRAM[62214] = 8'b10001011;
DRAM[62215] = 8'b10010000;
DRAM[62216] = 8'b10011001;
DRAM[62217] = 8'b10110100;
DRAM[62218] = 8'b11010100;
DRAM[62219] = 8'b11100111;
DRAM[62220] = 8'b11101110;
DRAM[62221] = 8'b11110001;
DRAM[62222] = 8'b11110010;
DRAM[62223] = 8'b11110001;
DRAM[62224] = 8'b11110010;
DRAM[62225] = 8'b11110000;
DRAM[62226] = 8'b11101111;
DRAM[62227] = 8'b11110000;
DRAM[62228] = 8'b11110011;
DRAM[62229] = 8'b11110100;
DRAM[62230] = 8'b11110000;
DRAM[62231] = 8'b11101100;
DRAM[62232] = 8'b11101000;
DRAM[62233] = 8'b11100001;
DRAM[62234] = 8'b11011011;
DRAM[62235] = 8'b11011100;
DRAM[62236] = 8'b11100000;
DRAM[62237] = 8'b11100001;
DRAM[62238] = 8'b11011011;
DRAM[62239] = 8'b11010101;
DRAM[62240] = 8'b11001101;
DRAM[62241] = 8'b11001011;
DRAM[62242] = 8'b11001001;
DRAM[62243] = 8'b11001010;
DRAM[62244] = 8'b11001101;
DRAM[62245] = 8'b11001101;
DRAM[62246] = 8'b11001010;
DRAM[62247] = 8'b11000111;
DRAM[62248] = 8'b11001010;
DRAM[62249] = 8'b10111110;
DRAM[62250] = 8'b10110011;
DRAM[62251] = 8'b10110001;
DRAM[62252] = 8'b10110110;
DRAM[62253] = 8'b10111001;
DRAM[62254] = 8'b10110100;
DRAM[62255] = 8'b10101101;
DRAM[62256] = 8'b10101100;
DRAM[62257] = 8'b10101001;
DRAM[62258] = 8'b10100011;
DRAM[62259] = 8'b10011011;
DRAM[62260] = 8'b10010100;
DRAM[62261] = 8'b10010011;
DRAM[62262] = 8'b10010111;
DRAM[62263] = 8'b10011011;
DRAM[62264] = 8'b10010111;
DRAM[62265] = 8'b10011010;
DRAM[62266] = 8'b10011111;
DRAM[62267] = 8'b10100010;
DRAM[62268] = 8'b10100100;
DRAM[62269] = 8'b10100000;
DRAM[62270] = 8'b10011001;
DRAM[62271] = 8'b10010010;
DRAM[62272] = 8'b10001010;
DRAM[62273] = 8'b10010000;
DRAM[62274] = 8'b10001111;
DRAM[62275] = 8'b10001000;
DRAM[62276] = 8'b10001000;
DRAM[62277] = 8'b10001101;
DRAM[62278] = 8'b10001010;
DRAM[62279] = 8'b10000001;
DRAM[62280] = 8'b1110111;
DRAM[62281] = 8'b1110010;
DRAM[62282] = 8'b1110101;
DRAM[62283] = 8'b10000010;
DRAM[62284] = 8'b10001101;
DRAM[62285] = 8'b10001110;
DRAM[62286] = 8'b10001101;
DRAM[62287] = 8'b10010000;
DRAM[62288] = 8'b10001001;
DRAM[62289] = 8'b10001010;
DRAM[62290] = 8'b1111001;
DRAM[62291] = 8'b10001010;
DRAM[62292] = 8'b10001011;
DRAM[62293] = 8'b1111010;
DRAM[62294] = 8'b10000110;
DRAM[62295] = 8'b10000000;
DRAM[62296] = 8'b10000100;
DRAM[62297] = 8'b1110101;
DRAM[62298] = 8'b1110011;
DRAM[62299] = 8'b1111111;
DRAM[62300] = 8'b10000001;
DRAM[62301] = 8'b1110101;
DRAM[62302] = 8'b1110001;
DRAM[62303] = 8'b1111010;
DRAM[62304] = 8'b1110100;
DRAM[62305] = 8'b1100110;
DRAM[62306] = 8'b1101011;
DRAM[62307] = 8'b1111010;
DRAM[62308] = 8'b1111001;
DRAM[62309] = 8'b1110100;
DRAM[62310] = 8'b1110100;
DRAM[62311] = 8'b1110011;
DRAM[62312] = 8'b1100101;
DRAM[62313] = 8'b10000000;
DRAM[62314] = 8'b10000101;
DRAM[62315] = 8'b1101100;
DRAM[62316] = 8'b1100000;
DRAM[62317] = 8'b1101100;
DRAM[62318] = 8'b1101111;
DRAM[62319] = 8'b1100011;
DRAM[62320] = 8'b1110001;
DRAM[62321] = 8'b1101111;
DRAM[62322] = 8'b1100111;
DRAM[62323] = 8'b1011110;
DRAM[62324] = 8'b1011110;
DRAM[62325] = 8'b1101010;
DRAM[62326] = 8'b1110100;
DRAM[62327] = 8'b1111001;
DRAM[62328] = 8'b1101010;
DRAM[62329] = 8'b1100111;
DRAM[62330] = 8'b1011110;
DRAM[62331] = 8'b1110000;
DRAM[62332] = 8'b1111001;
DRAM[62333] = 8'b1110000;
DRAM[62334] = 8'b1110010;
DRAM[62335] = 8'b1101001;
DRAM[62336] = 8'b1101100;
DRAM[62337] = 8'b1110000;
DRAM[62338] = 8'b1110011;
DRAM[62339] = 8'b1110001;
DRAM[62340] = 8'b1101101;
DRAM[62341] = 8'b1101100;
DRAM[62342] = 8'b1101111;
DRAM[62343] = 8'b1110010;
DRAM[62344] = 8'b1101101;
DRAM[62345] = 8'b1101010;
DRAM[62346] = 8'b1100110;
DRAM[62347] = 8'b1100100;
DRAM[62348] = 8'b1100111;
DRAM[62349] = 8'b1101011;
DRAM[62350] = 8'b1101001;
DRAM[62351] = 8'b1100011;
DRAM[62352] = 8'b1101010;
DRAM[62353] = 8'b1101011;
DRAM[62354] = 8'b1100111;
DRAM[62355] = 8'b1100111;
DRAM[62356] = 8'b1101100;
DRAM[62357] = 8'b1100110;
DRAM[62358] = 8'b1100100;
DRAM[62359] = 8'b1110000;
DRAM[62360] = 8'b1101001;
DRAM[62361] = 8'b1101110;
DRAM[62362] = 8'b1101110;
DRAM[62363] = 8'b1100111;
DRAM[62364] = 8'b1100101;
DRAM[62365] = 8'b1101011;
DRAM[62366] = 8'b1110101;
DRAM[62367] = 8'b1111011;
DRAM[62368] = 8'b1111001;
DRAM[62369] = 8'b1111110;
DRAM[62370] = 8'b10000010;
DRAM[62371] = 8'b10000011;
DRAM[62372] = 8'b1111111;
DRAM[62373] = 8'b1111101;
DRAM[62374] = 8'b1111110;
DRAM[62375] = 8'b10000000;
DRAM[62376] = 8'b10000110;
DRAM[62377] = 8'b10000111;
DRAM[62378] = 8'b10010000;
DRAM[62379] = 8'b10011011;
DRAM[62380] = 8'b10011001;
DRAM[62381] = 8'b10010001;
DRAM[62382] = 8'b10010010;
DRAM[62383] = 8'b10011011;
DRAM[62384] = 8'b10101001;
DRAM[62385] = 8'b10101010;
DRAM[62386] = 8'b10101100;
DRAM[62387] = 8'b10101110;
DRAM[62388] = 8'b10110010;
DRAM[62389] = 8'b10110110;
DRAM[62390] = 8'b10111011;
DRAM[62391] = 8'b10111110;
DRAM[62392] = 8'b11000100;
DRAM[62393] = 8'b11000110;
DRAM[62394] = 8'b11001001;
DRAM[62395] = 8'b11001010;
DRAM[62396] = 8'b11001100;
DRAM[62397] = 8'b11010001;
DRAM[62398] = 8'b11010111;
DRAM[62399] = 8'b11011010;
DRAM[62400] = 8'b11110010;
DRAM[62401] = 8'b11101101;
DRAM[62402] = 8'b11011010;
DRAM[62403] = 8'b11000000;
DRAM[62404] = 8'b10101110;
DRAM[62405] = 8'b10100101;
DRAM[62406] = 8'b10011010;
DRAM[62407] = 8'b10001110;
DRAM[62408] = 8'b10010011;
DRAM[62409] = 8'b10001111;
DRAM[62410] = 8'b10001011;
DRAM[62411] = 8'b10001000;
DRAM[62412] = 8'b10000101;
DRAM[62413] = 8'b10000001;
DRAM[62414] = 8'b1111101;
DRAM[62415] = 8'b1111010;
DRAM[62416] = 8'b1110110;
DRAM[62417] = 8'b1110101;
DRAM[62418] = 8'b1110100;
DRAM[62419] = 8'b1110010;
DRAM[62420] = 8'b1101111;
DRAM[62421] = 8'b1101100;
DRAM[62422] = 8'b1101001;
DRAM[62423] = 8'b1100111;
DRAM[62424] = 8'b1101000;
DRAM[62425] = 8'b1101000;
DRAM[62426] = 8'b1101000;
DRAM[62427] = 8'b1101000;
DRAM[62428] = 8'b1101000;
DRAM[62429] = 8'b1101001;
DRAM[62430] = 8'b1101001;
DRAM[62431] = 8'b1101001;
DRAM[62432] = 8'b1100101;
DRAM[62433] = 8'b1100110;
DRAM[62434] = 8'b1100110;
DRAM[62435] = 8'b1100110;
DRAM[62436] = 8'b1100110;
DRAM[62437] = 8'b1100111;
DRAM[62438] = 8'b1100111;
DRAM[62439] = 8'b1100111;
DRAM[62440] = 8'b1101001;
DRAM[62441] = 8'b1101000;
DRAM[62442] = 8'b1101000;
DRAM[62443] = 8'b1100111;
DRAM[62444] = 8'b1100111;
DRAM[62445] = 8'b1101000;
DRAM[62446] = 8'b1101000;
DRAM[62447] = 8'b1101001;
DRAM[62448] = 8'b1101010;
DRAM[62449] = 8'b1101011;
DRAM[62450] = 8'b1101110;
DRAM[62451] = 8'b1110000;
DRAM[62452] = 8'b1110001;
DRAM[62453] = 8'b1110000;
DRAM[62454] = 8'b1101111;
DRAM[62455] = 8'b1101110;
DRAM[62456] = 8'b1101010;
DRAM[62457] = 8'b1101001;
DRAM[62458] = 8'b1101001;
DRAM[62459] = 8'b1100111;
DRAM[62460] = 8'b1100110;
DRAM[62461] = 8'b1100101;
DRAM[62462] = 8'b1100100;
DRAM[62463] = 8'b1100100;
DRAM[62464] = 8'b10010001;
DRAM[62465] = 8'b10001100;
DRAM[62466] = 8'b10001010;
DRAM[62467] = 8'b10001011;
DRAM[62468] = 8'b10001010;
DRAM[62469] = 8'b10001001;
DRAM[62470] = 8'b10001111;
DRAM[62471] = 8'b10011000;
DRAM[62472] = 8'b10101101;
DRAM[62473] = 8'b11000011;
DRAM[62474] = 8'b11011100;
DRAM[62475] = 8'b11101100;
DRAM[62476] = 8'b11110011;
DRAM[62477] = 8'b11110110;
DRAM[62478] = 8'b11110101;
DRAM[62479] = 8'b11110010;
DRAM[62480] = 8'b11110000;
DRAM[62481] = 8'b11101110;
DRAM[62482] = 8'b11101110;
DRAM[62483] = 8'b11110000;
DRAM[62484] = 8'b11110011;
DRAM[62485] = 8'b11110011;
DRAM[62486] = 8'b11101111;
DRAM[62487] = 8'b11101011;
DRAM[62488] = 8'b11100101;
DRAM[62489] = 8'b11011110;
DRAM[62490] = 8'b11010111;
DRAM[62491] = 8'b11010110;
DRAM[62492] = 8'b11011001;
DRAM[62493] = 8'b11011001;
DRAM[62494] = 8'b11010010;
DRAM[62495] = 8'b11001011;
DRAM[62496] = 8'b11001000;
DRAM[62497] = 8'b11001000;
DRAM[62498] = 8'b11000111;
DRAM[62499] = 8'b11000110;
DRAM[62500] = 8'b11000101;
DRAM[62501] = 8'b11000011;
DRAM[62502] = 8'b11000001;
DRAM[62503] = 8'b11000000;
DRAM[62504] = 8'b11000010;
DRAM[62505] = 8'b10111010;
DRAM[62506] = 8'b10110011;
DRAM[62507] = 8'b10110101;
DRAM[62508] = 8'b10111100;
DRAM[62509] = 8'b10111101;
DRAM[62510] = 8'b10110110;
DRAM[62511] = 8'b10101101;
DRAM[62512] = 8'b10111100;
DRAM[62513] = 8'b10110101;
DRAM[62514] = 8'b10101101;
DRAM[62515] = 8'b10100110;
DRAM[62516] = 8'b10100010;
DRAM[62517] = 8'b10100000;
DRAM[62518] = 8'b10011101;
DRAM[62519] = 8'b10011010;
DRAM[62520] = 8'b10011010;
DRAM[62521] = 8'b10011001;
DRAM[62522] = 8'b10011001;
DRAM[62523] = 8'b10011010;
DRAM[62524] = 8'b10011010;
DRAM[62525] = 8'b10010110;
DRAM[62526] = 8'b10010010;
DRAM[62527] = 8'b10001111;
DRAM[62528] = 8'b10001011;
DRAM[62529] = 8'b10010000;
DRAM[62530] = 8'b10001110;
DRAM[62531] = 8'b10001000;
DRAM[62532] = 8'b10001000;
DRAM[62533] = 8'b10001111;
DRAM[62534] = 8'b10001100;
DRAM[62535] = 8'b10000100;
DRAM[62536] = 8'b1110101;
DRAM[62537] = 8'b1110100;
DRAM[62538] = 8'b1110000;
DRAM[62539] = 8'b1110010;
DRAM[62540] = 8'b1111110;
DRAM[62541] = 8'b10001100;
DRAM[62542] = 8'b10001100;
DRAM[62543] = 8'b10000011;
DRAM[62544] = 8'b10010101;
DRAM[62545] = 8'b10010010;
DRAM[62546] = 8'b1111010;
DRAM[62547] = 8'b10000110;
DRAM[62548] = 8'b10000101;
DRAM[62549] = 8'b1110011;
DRAM[62550] = 8'b1111111;
DRAM[62551] = 8'b1111000;
DRAM[62552] = 8'b1111010;
DRAM[62553] = 8'b1111010;
DRAM[62554] = 8'b1111011;
DRAM[62555] = 8'b1111100;
DRAM[62556] = 8'b1111001;
DRAM[62557] = 8'b1110101;
DRAM[62558] = 8'b1110101;
DRAM[62559] = 8'b1110110;
DRAM[62560] = 8'b1110000;
DRAM[62561] = 8'b1011110;
DRAM[62562] = 8'b1100011;
DRAM[62563] = 8'b1111000;
DRAM[62564] = 8'b1111110;
DRAM[62565] = 8'b1111100;
DRAM[62566] = 8'b1111000;
DRAM[62567] = 8'b1110001;
DRAM[62568] = 8'b1100111;
DRAM[62569] = 8'b1101100;
DRAM[62570] = 8'b1110111;
DRAM[62571] = 8'b1111100;
DRAM[62572] = 8'b1110011;
DRAM[62573] = 8'b1100100;
DRAM[62574] = 8'b1100010;
DRAM[62575] = 8'b1101010;
DRAM[62576] = 8'b1111000;
DRAM[62577] = 8'b1110001;
DRAM[62578] = 8'b1100100;
DRAM[62579] = 8'b1011010;
DRAM[62580] = 8'b1011011;
DRAM[62581] = 8'b1100100;
DRAM[62582] = 8'b1101000;
DRAM[62583] = 8'b1100110;
DRAM[62584] = 8'b1101111;
DRAM[62585] = 8'b1110010;
DRAM[62586] = 8'b1100010;
DRAM[62587] = 8'b1100101;
DRAM[62588] = 8'b1101110;
DRAM[62589] = 8'b1110101;
DRAM[62590] = 8'b1111111;
DRAM[62591] = 8'b1110001;
DRAM[62592] = 8'b1100101;
DRAM[62593] = 8'b1100011;
DRAM[62594] = 8'b1100100;
DRAM[62595] = 8'b1101011;
DRAM[62596] = 8'b1110011;
DRAM[62597] = 8'b1110110;
DRAM[62598] = 8'b1110101;
DRAM[62599] = 8'b1110011;
DRAM[62600] = 8'b1110011;
DRAM[62601] = 8'b1110000;
DRAM[62602] = 8'b1101001;
DRAM[62603] = 8'b1100011;
DRAM[62604] = 8'b1100101;
DRAM[62605] = 8'b1101001;
DRAM[62606] = 8'b1100101;
DRAM[62607] = 8'b1011100;
DRAM[62608] = 8'b1101110;
DRAM[62609] = 8'b1101100;
DRAM[62610] = 8'b1100101;
DRAM[62611] = 8'b1100111;
DRAM[62612] = 8'b1110001;
DRAM[62613] = 8'b1101110;
DRAM[62614] = 8'b1100111;
DRAM[62615] = 8'b1101011;
DRAM[62616] = 8'b1101010;
DRAM[62617] = 8'b1101101;
DRAM[62618] = 8'b1101110;
DRAM[62619] = 8'b1101011;
DRAM[62620] = 8'b1101100;
DRAM[62621] = 8'b1110010;
DRAM[62622] = 8'b1110111;
DRAM[62623] = 8'b1111000;
DRAM[62624] = 8'b1111001;
DRAM[62625] = 8'b1111110;
DRAM[62626] = 8'b10000010;
DRAM[62627] = 8'b10000011;
DRAM[62628] = 8'b10000001;
DRAM[62629] = 8'b1111111;
DRAM[62630] = 8'b1111110;
DRAM[62631] = 8'b1111111;
DRAM[62632] = 8'b10001000;
DRAM[62633] = 8'b10000011;
DRAM[62634] = 8'b10000110;
DRAM[62635] = 8'b10010010;
DRAM[62636] = 8'b10011000;
DRAM[62637] = 8'b10010100;
DRAM[62638] = 8'b10010100;
DRAM[62639] = 8'b10011010;
DRAM[62640] = 8'b10011100;
DRAM[62641] = 8'b10100011;
DRAM[62642] = 8'b10101010;
DRAM[62643] = 8'b10101100;
DRAM[62644] = 8'b10101011;
DRAM[62645] = 8'b10101101;
DRAM[62646] = 8'b10110101;
DRAM[62647] = 8'b10111011;
DRAM[62648] = 8'b10111100;
DRAM[62649] = 8'b10111110;
DRAM[62650] = 8'b11000010;
DRAM[62651] = 8'b11001000;
DRAM[62652] = 8'b11001110;
DRAM[62653] = 8'b11010101;
DRAM[62654] = 8'b11011101;
DRAM[62655] = 8'b11100100;
DRAM[62656] = 8'b11101011;
DRAM[62657] = 8'b11101010;
DRAM[62658] = 8'b11011010;
DRAM[62659] = 8'b10111111;
DRAM[62660] = 8'b10101010;
DRAM[62661] = 8'b10011110;
DRAM[62662] = 8'b10010100;
DRAM[62663] = 8'b10001010;
DRAM[62664] = 8'b10010000;
DRAM[62665] = 8'b10001101;
DRAM[62666] = 8'b10001000;
DRAM[62667] = 8'b10000101;
DRAM[62668] = 8'b10000010;
DRAM[62669] = 8'b1111111;
DRAM[62670] = 8'b1111010;
DRAM[62671] = 8'b1110111;
DRAM[62672] = 8'b1110011;
DRAM[62673] = 8'b1110011;
DRAM[62674] = 8'b1110001;
DRAM[62675] = 8'b1101111;
DRAM[62676] = 8'b1101100;
DRAM[62677] = 8'b1101001;
DRAM[62678] = 8'b1100110;
DRAM[62679] = 8'b1100101;
DRAM[62680] = 8'b1100100;
DRAM[62681] = 8'b1100100;
DRAM[62682] = 8'b1100101;
DRAM[62683] = 8'b1100101;
DRAM[62684] = 8'b1100110;
DRAM[62685] = 8'b1100111;
DRAM[62686] = 8'b1100111;
DRAM[62687] = 8'b1100111;
DRAM[62688] = 8'b1100100;
DRAM[62689] = 8'b1100101;
DRAM[62690] = 8'b1100101;
DRAM[62691] = 8'b1100110;
DRAM[62692] = 8'b1100110;
DRAM[62693] = 8'b1100111;
DRAM[62694] = 8'b1100111;
DRAM[62695] = 8'b1100111;
DRAM[62696] = 8'b1101001;
DRAM[62697] = 8'b1101000;
DRAM[62698] = 8'b1101000;
DRAM[62699] = 8'b1100111;
DRAM[62700] = 8'b1100111;
DRAM[62701] = 8'b1101000;
DRAM[62702] = 8'b1101000;
DRAM[62703] = 8'b1101001;
DRAM[62704] = 8'b1101001;
DRAM[62705] = 8'b1101011;
DRAM[62706] = 8'b1101110;
DRAM[62707] = 8'b1110000;
DRAM[62708] = 8'b1110001;
DRAM[62709] = 8'b1110000;
DRAM[62710] = 8'b1101111;
DRAM[62711] = 8'b1101101;
DRAM[62712] = 8'b1101010;
DRAM[62713] = 8'b1101001;
DRAM[62714] = 8'b1101001;
DRAM[62715] = 8'b1100111;
DRAM[62716] = 8'b1100110;
DRAM[62717] = 8'b1100101;
DRAM[62718] = 8'b1100100;
DRAM[62719] = 8'b1100100;
DRAM[62720] = 8'b10010010;
DRAM[62721] = 8'b10001100;
DRAM[62722] = 8'b10001010;
DRAM[62723] = 8'b10001100;
DRAM[62724] = 8'b10001011;
DRAM[62725] = 8'b10001011;
DRAM[62726] = 8'b10010100;
DRAM[62727] = 8'b10100001;
DRAM[62728] = 8'b10111101;
DRAM[62729] = 8'b11001110;
DRAM[62730] = 8'b11100010;
DRAM[62731] = 8'b11101110;
DRAM[62732] = 8'b11110100;
DRAM[62733] = 8'b11110111;
DRAM[62734] = 8'b11110101;
DRAM[62735] = 8'b11110001;
DRAM[62736] = 8'b11101111;
DRAM[62737] = 8'b11101110;
DRAM[62738] = 8'b11101101;
DRAM[62739] = 8'b11101111;
DRAM[62740] = 8'b11110010;
DRAM[62741] = 8'b11110001;
DRAM[62742] = 8'b11101101;
DRAM[62743] = 8'b11101000;
DRAM[62744] = 8'b11100101;
DRAM[62745] = 8'b11011111;
DRAM[62746] = 8'b11011000;
DRAM[62747] = 8'b11010110;
DRAM[62748] = 8'b11010110;
DRAM[62749] = 8'b11010011;
DRAM[62750] = 8'b11001101;
DRAM[62751] = 8'b11000111;
DRAM[62752] = 8'b11001001;
DRAM[62753] = 8'b11001001;
DRAM[62754] = 8'b11001000;
DRAM[62755] = 8'b11000101;
DRAM[62756] = 8'b11000001;
DRAM[62757] = 8'b10111110;
DRAM[62758] = 8'b10111110;
DRAM[62759] = 8'b10111110;
DRAM[62760] = 8'b10110110;
DRAM[62761] = 8'b10111011;
DRAM[62762] = 8'b10111111;
DRAM[62763] = 8'b11000001;
DRAM[62764] = 8'b10111111;
DRAM[62765] = 8'b10111100;
DRAM[62766] = 8'b10111011;
DRAM[62767] = 8'b10111011;
DRAM[62768] = 8'b10110110;
DRAM[62769] = 8'b10110011;
DRAM[62770] = 8'b10110001;
DRAM[62771] = 8'b10110001;
DRAM[62772] = 8'b10110010;
DRAM[62773] = 8'b10101101;
DRAM[62774] = 8'b10100101;
DRAM[62775] = 8'b10011101;
DRAM[62776] = 8'b10100011;
DRAM[62777] = 8'b10011011;
DRAM[62778] = 8'b10010011;
DRAM[62779] = 8'b10001110;
DRAM[62780] = 8'b10001011;
DRAM[62781] = 8'b10001010;
DRAM[62782] = 8'b10001110;
DRAM[62783] = 8'b10010101;
DRAM[62784] = 8'b10001011;
DRAM[62785] = 8'b10001110;
DRAM[62786] = 8'b10001110;
DRAM[62787] = 8'b10001011;
DRAM[62788] = 8'b10001011;
DRAM[62789] = 8'b10001101;
DRAM[62790] = 8'b10001101;
DRAM[62791] = 8'b10001011;
DRAM[62792] = 8'b1111001;
DRAM[62793] = 8'b1111110;
DRAM[62794] = 8'b1111010;
DRAM[62795] = 8'b1110010;
DRAM[62796] = 8'b1111000;
DRAM[62797] = 8'b10001000;
DRAM[62798] = 8'b10001011;
DRAM[62799] = 8'b10000011;
DRAM[62800] = 8'b10001111;
DRAM[62801] = 8'b10001010;
DRAM[62802] = 8'b1111100;
DRAM[62803] = 8'b1111111;
DRAM[62804] = 8'b1111111;
DRAM[62805] = 8'b1111001;
DRAM[62806] = 8'b1111110;
DRAM[62807] = 8'b1111011;
DRAM[62808] = 8'b1110110;
DRAM[62809] = 8'b1111000;
DRAM[62810] = 8'b1110110;
DRAM[62811] = 8'b1110100;
DRAM[62812] = 8'b1111010;
DRAM[62813] = 8'b10000010;
DRAM[62814] = 8'b1111100;
DRAM[62815] = 8'b1101110;
DRAM[62816] = 8'b1101010;
DRAM[62817] = 8'b1101000;
DRAM[62818] = 8'b1101011;
DRAM[62819] = 8'b1101110;
DRAM[62820] = 8'b1110110;
DRAM[62821] = 8'b10000100;
DRAM[62822] = 8'b10000000;
DRAM[62823] = 8'b1100111;
DRAM[62824] = 8'b1101101;
DRAM[62825] = 8'b1101001;
DRAM[62826] = 8'b1100110;
DRAM[62827] = 8'b1101000;
DRAM[62828] = 8'b1101101;
DRAM[62829] = 8'b1101111;
DRAM[62830] = 8'b1101101;
DRAM[62831] = 8'b1101011;
DRAM[62832] = 8'b1100001;
DRAM[62833] = 8'b1100111;
DRAM[62834] = 8'b1101101;
DRAM[62835] = 8'b1101011;
DRAM[62836] = 8'b1100101;
DRAM[62837] = 8'b1100010;
DRAM[62838] = 8'b1100101;
DRAM[62839] = 8'b1101011;
DRAM[62840] = 8'b1101010;
DRAM[62841] = 8'b1111010;
DRAM[62842] = 8'b1110000;
DRAM[62843] = 8'b1101001;
DRAM[62844] = 8'b1100101;
DRAM[62845] = 8'b1101101;
DRAM[62846] = 8'b10000010;
DRAM[62847] = 8'b1111110;
DRAM[62848] = 8'b1101000;
DRAM[62849] = 8'b1011111;
DRAM[62850] = 8'b1011100;
DRAM[62851] = 8'b1100110;
DRAM[62852] = 8'b1110011;
DRAM[62853] = 8'b1111000;
DRAM[62854] = 8'b1110100;
DRAM[62855] = 8'b1110000;
DRAM[62856] = 8'b1110110;
DRAM[62857] = 8'b1110100;
DRAM[62858] = 8'b1101100;
DRAM[62859] = 8'b1100100;
DRAM[62860] = 8'b1100100;
DRAM[62861] = 8'b1101001;
DRAM[62862] = 8'b1100101;
DRAM[62863] = 8'b1011100;
DRAM[62864] = 8'b1101100;
DRAM[62865] = 8'b1101110;
DRAM[62866] = 8'b1100110;
DRAM[62867] = 8'b1100100;
DRAM[62868] = 8'b1110001;
DRAM[62869] = 8'b1110100;
DRAM[62870] = 8'b1101010;
DRAM[62871] = 8'b1100101;
DRAM[62872] = 8'b1101101;
DRAM[62873] = 8'b1110001;
DRAM[62874] = 8'b1110011;
DRAM[62875] = 8'b1110010;
DRAM[62876] = 8'b1110100;
DRAM[62877] = 8'b1111001;
DRAM[62878] = 8'b1111011;
DRAM[62879] = 8'b1111001;
DRAM[62880] = 8'b1111011;
DRAM[62881] = 8'b1111110;
DRAM[62882] = 8'b10000001;
DRAM[62883] = 8'b10000011;
DRAM[62884] = 8'b10000001;
DRAM[62885] = 8'b10000000;
DRAM[62886] = 8'b1111111;
DRAM[62887] = 8'b1111111;
DRAM[62888] = 8'b10001000;
DRAM[62889] = 8'b10000011;
DRAM[62890] = 8'b10000011;
DRAM[62891] = 8'b10001100;
DRAM[62892] = 8'b10010101;
DRAM[62893] = 8'b10011000;
DRAM[62894] = 8'b10011001;
DRAM[62895] = 8'b10011010;
DRAM[62896] = 8'b10010010;
DRAM[62897] = 8'b10011001;
DRAM[62898] = 8'b10100010;
DRAM[62899] = 8'b10100110;
DRAM[62900] = 8'b10100111;
DRAM[62901] = 8'b10101100;
DRAM[62902] = 8'b10110101;
DRAM[62903] = 8'b10111100;
DRAM[62904] = 8'b10111010;
DRAM[62905] = 8'b10111001;
DRAM[62906] = 8'b10111101;
DRAM[62907] = 8'b11000100;
DRAM[62908] = 8'b11001011;
DRAM[62909] = 8'b11010001;
DRAM[62910] = 8'b11011100;
DRAM[62911] = 8'b11100110;
DRAM[62912] = 8'b11100100;
DRAM[62913] = 8'b11100111;
DRAM[62914] = 8'b11011110;
DRAM[62915] = 8'b11001000;
DRAM[62916] = 8'b10110100;
DRAM[62917] = 8'b10101000;
DRAM[62918] = 8'b10011100;
DRAM[62919] = 8'b10010000;
DRAM[62920] = 8'b10010000;
DRAM[62921] = 8'b10001100;
DRAM[62922] = 8'b10000111;
DRAM[62923] = 8'b10000011;
DRAM[62924] = 8'b1111111;
DRAM[62925] = 8'b1111010;
DRAM[62926] = 8'b1110101;
DRAM[62927] = 8'b1110010;
DRAM[62928] = 8'b1110000;
DRAM[62929] = 8'b1101111;
DRAM[62930] = 8'b1101110;
DRAM[62931] = 8'b1101100;
DRAM[62932] = 8'b1101001;
DRAM[62933] = 8'b1100110;
DRAM[62934] = 8'b1100011;
DRAM[62935] = 8'b1100001;
DRAM[62936] = 8'b1100001;
DRAM[62937] = 8'b1100001;
DRAM[62938] = 8'b1100010;
DRAM[62939] = 8'b1100011;
DRAM[62940] = 8'b1100100;
DRAM[62941] = 8'b1100101;
DRAM[62942] = 8'b1100110;
DRAM[62943] = 8'b1100110;
DRAM[62944] = 8'b1100100;
DRAM[62945] = 8'b1100100;
DRAM[62946] = 8'b1100100;
DRAM[62947] = 8'b1100101;
DRAM[62948] = 8'b1100110;
DRAM[62949] = 8'b1100110;
DRAM[62950] = 8'b1100111;
DRAM[62951] = 8'b1100111;
DRAM[62952] = 8'b1101001;
DRAM[62953] = 8'b1101000;
DRAM[62954] = 8'b1101000;
DRAM[62955] = 8'b1100111;
DRAM[62956] = 8'b1100111;
DRAM[62957] = 8'b1101000;
DRAM[62958] = 8'b1101000;
DRAM[62959] = 8'b1101001;
DRAM[62960] = 8'b1101001;
DRAM[62961] = 8'b1101011;
DRAM[62962] = 8'b1101101;
DRAM[62963] = 8'b1101111;
DRAM[62964] = 8'b1110000;
DRAM[62965] = 8'b1110000;
DRAM[62966] = 8'b1101110;
DRAM[62967] = 8'b1101101;
DRAM[62968] = 8'b1101011;
DRAM[62969] = 8'b1101010;
DRAM[62970] = 8'b1101001;
DRAM[62971] = 8'b1101000;
DRAM[62972] = 8'b1100111;
DRAM[62973] = 8'b1100110;
DRAM[62974] = 8'b1100101;
DRAM[62975] = 8'b1100100;
DRAM[62976] = 8'b10010010;
DRAM[62977] = 8'b10001100;
DRAM[62978] = 8'b10001010;
DRAM[62979] = 8'b10001110;
DRAM[62980] = 8'b10001110;
DRAM[62981] = 8'b10001101;
DRAM[62982] = 8'b10011001;
DRAM[62983] = 8'b10101010;
DRAM[62984] = 8'b11000011;
DRAM[62985] = 8'b11010101;
DRAM[62986] = 8'b11101000;
DRAM[62987] = 8'b11110000;
DRAM[62988] = 8'b11110010;
DRAM[62989] = 8'b11110011;
DRAM[62990] = 8'b11110010;
DRAM[62991] = 8'b11110000;
DRAM[62992] = 8'b11101111;
DRAM[62993] = 8'b11101110;
DRAM[62994] = 8'b11101101;
DRAM[62995] = 8'b11101111;
DRAM[62996] = 8'b11110001;
DRAM[62997] = 8'b11110000;
DRAM[62998] = 8'b11101010;
DRAM[62999] = 8'b11100101;
DRAM[63000] = 8'b11100010;
DRAM[63001] = 8'b11011110;
DRAM[63002] = 8'b11011010;
DRAM[63003] = 8'b11010110;
DRAM[63004] = 8'b11010011;
DRAM[63005] = 8'b11001111;
DRAM[63006] = 8'b11001011;
DRAM[63007] = 8'b11000111;
DRAM[63008] = 8'b10111111;
DRAM[63009] = 8'b11000000;
DRAM[63010] = 8'b10111111;
DRAM[63011] = 8'b10111010;
DRAM[63012] = 8'b10110101;
DRAM[63013] = 8'b10110010;
DRAM[63014] = 8'b10110100;
DRAM[63015] = 8'b10110111;
DRAM[63016] = 8'b10101110;
DRAM[63017] = 8'b10110010;
DRAM[63018] = 8'b10110111;
DRAM[63019] = 8'b10110111;
DRAM[63020] = 8'b10110100;
DRAM[63021] = 8'b10101111;
DRAM[63022] = 8'b10101101;
DRAM[63023] = 8'b10101101;
DRAM[63024] = 8'b10100000;
DRAM[63025] = 8'b10011111;
DRAM[63026] = 8'b10100000;
DRAM[63027] = 8'b10100000;
DRAM[63028] = 8'b10011111;
DRAM[63029] = 8'b10011101;
DRAM[63030] = 8'b10011010;
DRAM[63031] = 8'b10011000;
DRAM[63032] = 8'b10011011;
DRAM[63033] = 8'b10010101;
DRAM[63034] = 8'b10001111;
DRAM[63035] = 8'b10001101;
DRAM[63036] = 8'b10001001;
DRAM[63037] = 8'b10001001;
DRAM[63038] = 8'b10010001;
DRAM[63039] = 8'b10011100;
DRAM[63040] = 8'b10010101;
DRAM[63041] = 8'b10010101;
DRAM[63042] = 8'b10010110;
DRAM[63043] = 8'b10010110;
DRAM[63044] = 8'b10010000;
DRAM[63045] = 8'b10000111;
DRAM[63046] = 8'b10000101;
DRAM[63047] = 8'b10001000;
DRAM[63048] = 8'b1111101;
DRAM[63049] = 8'b10000101;
DRAM[63050] = 8'b10001000;
DRAM[63051] = 8'b10000000;
DRAM[63052] = 8'b1110111;
DRAM[63053] = 8'b1110111;
DRAM[63054] = 8'b1111111;
DRAM[63055] = 8'b10000110;
DRAM[63056] = 8'b1111111;
DRAM[63057] = 8'b1111100;
DRAM[63058] = 8'b10000010;
DRAM[63059] = 8'b1111011;
DRAM[63060] = 8'b1111101;
DRAM[63061] = 8'b10000110;
DRAM[63062] = 8'b10000001;
DRAM[63063] = 8'b10000010;
DRAM[63064] = 8'b1110101;
DRAM[63065] = 8'b1110110;
DRAM[63066] = 8'b1110101;
DRAM[63067] = 8'b1110110;
DRAM[63068] = 8'b1111101;
DRAM[63069] = 8'b10000010;
DRAM[63070] = 8'b1111010;
DRAM[63071] = 8'b1101100;
DRAM[63072] = 8'b1101100;
DRAM[63073] = 8'b1101100;
DRAM[63074] = 8'b1110000;
DRAM[63075] = 8'b1101110;
DRAM[63076] = 8'b1110000;
DRAM[63077] = 8'b1111111;
DRAM[63078] = 8'b10000001;
DRAM[63079] = 8'b1101111;
DRAM[63080] = 8'b1110100;
DRAM[63081] = 8'b1110110;
DRAM[63082] = 8'b1101010;
DRAM[63083] = 8'b1011011;
DRAM[63084] = 8'b1100000;
DRAM[63085] = 8'b1110011;
DRAM[63086] = 8'b1111000;
DRAM[63087] = 8'b1101111;
DRAM[63088] = 8'b1010111;
DRAM[63089] = 8'b1100001;
DRAM[63090] = 8'b1110010;
DRAM[63091] = 8'b1111011;
DRAM[63092] = 8'b1110011;
DRAM[63093] = 8'b1101000;
DRAM[63094] = 8'b1101100;
DRAM[63095] = 8'b1111000;
DRAM[63096] = 8'b1101001;
DRAM[63097] = 8'b1110111;
DRAM[63098] = 8'b1110010;
DRAM[63099] = 8'b1110001;
DRAM[63100] = 8'b1101000;
DRAM[63101] = 8'b1100010;
DRAM[63102] = 8'b1110001;
DRAM[63103] = 8'b1110010;
DRAM[63104] = 8'b1110011;
DRAM[63105] = 8'b1100111;
DRAM[63106] = 8'b1011111;
DRAM[63107] = 8'b1100100;
DRAM[63108] = 8'b1101101;
DRAM[63109] = 8'b1101111;
DRAM[63110] = 8'b1101110;
DRAM[63111] = 8'b1101101;
DRAM[63112] = 8'b1110010;
DRAM[63113] = 8'b1110100;
DRAM[63114] = 8'b1101110;
DRAM[63115] = 8'b1100100;
DRAM[63116] = 8'b1100101;
DRAM[63117] = 8'b1101100;
DRAM[63118] = 8'b1101011;
DRAM[63119] = 8'b1100011;
DRAM[63120] = 8'b1100111;
DRAM[63121] = 8'b1110011;
DRAM[63122] = 8'b1101101;
DRAM[63123] = 8'b1100100;
DRAM[63124] = 8'b1101110;
DRAM[63125] = 8'b1110110;
DRAM[63126] = 8'b1101101;
DRAM[63127] = 8'b1100100;
DRAM[63128] = 8'b1101100;
DRAM[63129] = 8'b1110100;
DRAM[63130] = 8'b1111001;
DRAM[63131] = 8'b1110110;
DRAM[63132] = 8'b1110011;
DRAM[63133] = 8'b1110110;
DRAM[63134] = 8'b1111011;
DRAM[63135] = 8'b1111101;
DRAM[63136] = 8'b1111101;
DRAM[63137] = 8'b1111111;
DRAM[63138] = 8'b10000001;
DRAM[63139] = 8'b10000010;
DRAM[63140] = 8'b10000001;
DRAM[63141] = 8'b10000000;
DRAM[63142] = 8'b10000000;
DRAM[63143] = 8'b10000000;
DRAM[63144] = 8'b10000100;
DRAM[63145] = 8'b10001000;
DRAM[63146] = 8'b10001010;
DRAM[63147] = 8'b10001101;
DRAM[63148] = 8'b10010011;
DRAM[63149] = 8'b10011010;
DRAM[63150] = 8'b10011100;
DRAM[63151] = 8'b10011001;
DRAM[63152] = 8'b10011000;
DRAM[63153] = 8'b10011000;
DRAM[63154] = 8'b10011001;
DRAM[63155] = 8'b10011011;
DRAM[63156] = 8'b10100001;
DRAM[63157] = 8'b10100111;
DRAM[63158] = 8'b10101100;
DRAM[63159] = 8'b10110000;
DRAM[63160] = 8'b10110110;
DRAM[63161] = 8'b10110100;
DRAM[63162] = 8'b10110110;
DRAM[63163] = 8'b10111101;
DRAM[63164] = 8'b11000100;
DRAM[63165] = 8'b11001011;
DRAM[63166] = 8'b11011000;
DRAM[63167] = 8'b11100100;
DRAM[63168] = 8'b11100111;
DRAM[63169] = 8'b11100100;
DRAM[63170] = 8'b11010100;
DRAM[63171] = 8'b10111101;
DRAM[63172] = 8'b10101101;
DRAM[63173] = 8'b10100101;
DRAM[63174] = 8'b10011001;
DRAM[63175] = 8'b10001100;
DRAM[63176] = 8'b10001100;
DRAM[63177] = 8'b10001000;
DRAM[63178] = 8'b10000100;
DRAM[63179] = 8'b10000000;
DRAM[63180] = 8'b1111100;
DRAM[63181] = 8'b1111000;
DRAM[63182] = 8'b1110011;
DRAM[63183] = 8'b1110000;
DRAM[63184] = 8'b1101101;
DRAM[63185] = 8'b1101100;
DRAM[63186] = 8'b1101011;
DRAM[63187] = 8'b1101001;
DRAM[63188] = 8'b1100110;
DRAM[63189] = 8'b1100011;
DRAM[63190] = 8'b1100000;
DRAM[63191] = 8'b1011110;
DRAM[63192] = 8'b1011110;
DRAM[63193] = 8'b1011111;
DRAM[63194] = 8'b1100000;
DRAM[63195] = 8'b1100001;
DRAM[63196] = 8'b1100010;
DRAM[63197] = 8'b1100100;
DRAM[63198] = 8'b1100101;
DRAM[63199] = 8'b1100101;
DRAM[63200] = 8'b1100011;
DRAM[63201] = 8'b1100011;
DRAM[63202] = 8'b1100100;
DRAM[63203] = 8'b1100101;
DRAM[63204] = 8'b1100110;
DRAM[63205] = 8'b1100110;
DRAM[63206] = 8'b1100111;
DRAM[63207] = 8'b1100111;
DRAM[63208] = 8'b1101001;
DRAM[63209] = 8'b1101000;
DRAM[63210] = 8'b1101000;
DRAM[63211] = 8'b1100111;
DRAM[63212] = 8'b1100111;
DRAM[63213] = 8'b1101000;
DRAM[63214] = 8'b1101000;
DRAM[63215] = 8'b1101001;
DRAM[63216] = 8'b1101001;
DRAM[63217] = 8'b1101010;
DRAM[63218] = 8'b1101101;
DRAM[63219] = 8'b1101111;
DRAM[63220] = 8'b1110000;
DRAM[63221] = 8'b1101111;
DRAM[63222] = 8'b1101110;
DRAM[63223] = 8'b1101101;
DRAM[63224] = 8'b1101100;
DRAM[63225] = 8'b1101011;
DRAM[63226] = 8'b1101010;
DRAM[63227] = 8'b1101001;
DRAM[63228] = 8'b1101000;
DRAM[63229] = 8'b1100111;
DRAM[63230] = 8'b1100110;
DRAM[63231] = 8'b1100101;
DRAM[63232] = 8'b10010011;
DRAM[63233] = 8'b10001100;
DRAM[63234] = 8'b10001011;
DRAM[63235] = 8'b10001111;
DRAM[63236] = 8'b10001111;
DRAM[63237] = 8'b10001111;
DRAM[63238] = 8'b10011101;
DRAM[63239] = 8'b10101111;
DRAM[63240] = 8'b11000110;
DRAM[63241] = 8'b11011011;
DRAM[63242] = 8'b11110000;
DRAM[63243] = 8'b11110111;
DRAM[63244] = 8'b11110100;
DRAM[63245] = 8'b11110010;
DRAM[63246] = 8'b11110010;
DRAM[63247] = 8'b11110011;
DRAM[63248] = 8'b11110000;
DRAM[63249] = 8'b11101110;
DRAM[63250] = 8'b11101110;
DRAM[63251] = 8'b11101111;
DRAM[63252] = 8'b11110001;
DRAM[63253] = 8'b11101111;
DRAM[63254] = 8'b11101001;
DRAM[63255] = 8'b11100100;
DRAM[63256] = 8'b11011001;
DRAM[63257] = 8'b11011000;
DRAM[63258] = 8'b11010101;
DRAM[63259] = 8'b11010001;
DRAM[63260] = 8'b11001100;
DRAM[63261] = 8'b11001000;
DRAM[63262] = 8'b11000101;
DRAM[63263] = 8'b11000011;
DRAM[63264] = 8'b11000110;
DRAM[63265] = 8'b11001000;
DRAM[63266] = 8'b11000111;
DRAM[63267] = 8'b11000010;
DRAM[63268] = 8'b10111100;
DRAM[63269] = 8'b10111010;
DRAM[63270] = 8'b10111101;
DRAM[63271] = 8'b11000001;
DRAM[63272] = 8'b11000011;
DRAM[63273] = 8'b10111011;
DRAM[63274] = 8'b10110100;
DRAM[63275] = 8'b10110110;
DRAM[63276] = 8'b10111010;
DRAM[63277] = 8'b10111000;
DRAM[63278] = 8'b10101101;
DRAM[63279] = 8'b10100010;
DRAM[63280] = 8'b10101111;
DRAM[63281] = 8'b10101101;
DRAM[63282] = 8'b10100111;
DRAM[63283] = 8'b10011110;
DRAM[63284] = 8'b10010110;
DRAM[63285] = 8'b10010101;
DRAM[63286] = 8'b10011010;
DRAM[63287] = 8'b10100000;
DRAM[63288] = 8'b10000001;
DRAM[63289] = 8'b10000001;
DRAM[63290] = 8'b10000110;
DRAM[63291] = 8'b10001011;
DRAM[63292] = 8'b10001010;
DRAM[63293] = 8'b10000111;
DRAM[63294] = 8'b10001110;
DRAM[63295] = 8'b10011001;
DRAM[63296] = 8'b10100110;
DRAM[63297] = 8'b10100010;
DRAM[63298] = 8'b10100001;
DRAM[63299] = 8'b10011110;
DRAM[63300] = 8'b10001110;
DRAM[63301] = 8'b1111000;
DRAM[63302] = 8'b1110000;
DRAM[63303] = 8'b1110100;
DRAM[63304] = 8'b1111100;
DRAM[63305] = 8'b10000011;
DRAM[63306] = 8'b10001100;
DRAM[63307] = 8'b10001000;
DRAM[63308] = 8'b1110001;
DRAM[63309] = 8'b1011111;
DRAM[63310] = 8'b1101010;
DRAM[63311] = 8'b10000001;
DRAM[63312] = 8'b1111101;
DRAM[63313] = 8'b1111011;
DRAM[63314] = 8'b10001100;
DRAM[63315] = 8'b1111100;
DRAM[63316] = 8'b1111011;
DRAM[63317] = 8'b10001011;
DRAM[63318] = 8'b1111010;
DRAM[63319] = 8'b1111101;
DRAM[63320] = 8'b1110011;
DRAM[63321] = 8'b1110111;
DRAM[63322] = 8'b1111100;
DRAM[63323] = 8'b1111111;
DRAM[63324] = 8'b1111100;
DRAM[63325] = 8'b1110101;
DRAM[63326] = 8'b1110001;
DRAM[63327] = 8'b1110000;
DRAM[63328] = 8'b1110100;
DRAM[63329] = 8'b1100110;
DRAM[63330] = 8'b1101011;
DRAM[63331] = 8'b1110111;
DRAM[63332] = 8'b1110100;
DRAM[63333] = 8'b1110010;
DRAM[63334] = 8'b1111100;
DRAM[63335] = 8'b10000011;
DRAM[63336] = 8'b1111001;
DRAM[63337] = 8'b1101111;
DRAM[63338] = 8'b1110010;
DRAM[63339] = 8'b1111100;
DRAM[63340] = 8'b1110101;
DRAM[63341] = 8'b1100010;
DRAM[63342] = 8'b1100101;
DRAM[63343] = 8'b1111000;
DRAM[63344] = 8'b1110100;
DRAM[63345] = 8'b1100100;
DRAM[63346] = 8'b1100010;
DRAM[63347] = 8'b1110100;
DRAM[63348] = 8'b1111111;
DRAM[63349] = 8'b1110110;
DRAM[63350] = 8'b1101010;
DRAM[63351] = 8'b1100110;
DRAM[63352] = 8'b1110001;
DRAM[63353] = 8'b1110000;
DRAM[63354] = 8'b1101000;
DRAM[63355] = 8'b1110101;
DRAM[63356] = 8'b1110001;
DRAM[63357] = 8'b1011100;
DRAM[63358] = 8'b1011100;
DRAM[63359] = 8'b1011000;
DRAM[63360] = 8'b1110110;
DRAM[63361] = 8'b1101001;
DRAM[63362] = 8'b1100000;
DRAM[63363] = 8'b1100010;
DRAM[63364] = 8'b1101000;
DRAM[63365] = 8'b1101011;
DRAM[63366] = 8'b1101111;
DRAM[63367] = 8'b1110100;
DRAM[63368] = 8'b1101101;
DRAM[63369] = 8'b1110010;
DRAM[63370] = 8'b1101110;
DRAM[63371] = 8'b1100101;
DRAM[63372] = 8'b1100110;
DRAM[63373] = 8'b1101111;
DRAM[63374] = 8'b1110001;
DRAM[63375] = 8'b1101010;
DRAM[63376] = 8'b1100100;
DRAM[63377] = 8'b1111000;
DRAM[63378] = 8'b1110101;
DRAM[63379] = 8'b1100110;
DRAM[63380] = 8'b1101101;
DRAM[63381] = 8'b1111000;
DRAM[63382] = 8'b1110001;
DRAM[63383] = 8'b1100110;
DRAM[63384] = 8'b1101001;
DRAM[63385] = 8'b1110100;
DRAM[63386] = 8'b1111011;
DRAM[63387] = 8'b1110101;
DRAM[63388] = 8'b1101110;
DRAM[63389] = 8'b1101111;
DRAM[63390] = 8'b1111000;
DRAM[63391] = 8'b1111111;
DRAM[63392] = 8'b1111110;
DRAM[63393] = 8'b1111111;
DRAM[63394] = 8'b10000000;
DRAM[63395] = 8'b10000001;
DRAM[63396] = 8'b10000001;
DRAM[63397] = 8'b10000001;
DRAM[63398] = 8'b10000001;
DRAM[63399] = 8'b10000001;
DRAM[63400] = 8'b10000001;
DRAM[63401] = 8'b10001100;
DRAM[63402] = 8'b10010011;
DRAM[63403] = 8'b10010000;
DRAM[63404] = 8'b10010010;
DRAM[63405] = 8'b10011010;
DRAM[63406] = 8'b10011101;
DRAM[63407] = 8'b10011001;
DRAM[63408] = 8'b10100011;
DRAM[63409] = 8'b10011001;
DRAM[63410] = 8'b10010000;
DRAM[63411] = 8'b10001110;
DRAM[63412] = 8'b10010101;
DRAM[63413] = 8'b10011011;
DRAM[63414] = 8'b10011011;
DRAM[63415] = 8'b10011001;
DRAM[63416] = 8'b10101000;
DRAM[63417] = 8'b10100110;
DRAM[63418] = 8'b10101010;
DRAM[63419] = 8'b10110110;
DRAM[63420] = 8'b11000001;
DRAM[63421] = 8'b11001100;
DRAM[63422] = 8'b11011101;
DRAM[63423] = 8'b11101100;
DRAM[63424] = 8'b11110001;
DRAM[63425] = 8'b11100010;
DRAM[63426] = 8'b11000100;
DRAM[63427] = 8'b10100110;
DRAM[63428] = 8'b10010111;
DRAM[63429] = 8'b10010011;
DRAM[63430] = 8'b10001011;
DRAM[63431] = 8'b1111110;
DRAM[63432] = 8'b10000101;
DRAM[63433] = 8'b10000010;
DRAM[63434] = 8'b1111111;
DRAM[63435] = 8'b1111101;
DRAM[63436] = 8'b1111011;
DRAM[63437] = 8'b1111001;
DRAM[63438] = 8'b1110101;
DRAM[63439] = 8'b1110011;
DRAM[63440] = 8'b1101011;
DRAM[63441] = 8'b1101010;
DRAM[63442] = 8'b1101001;
DRAM[63443] = 8'b1100111;
DRAM[63444] = 8'b1100100;
DRAM[63445] = 8'b1100001;
DRAM[63446] = 8'b1011110;
DRAM[63447] = 8'b1011100;
DRAM[63448] = 8'b1011101;
DRAM[63449] = 8'b1011101;
DRAM[63450] = 8'b1011111;
DRAM[63451] = 8'b1100000;
DRAM[63452] = 8'b1100010;
DRAM[63453] = 8'b1100011;
DRAM[63454] = 8'b1100100;
DRAM[63455] = 8'b1100101;
DRAM[63456] = 8'b1100010;
DRAM[63457] = 8'b1100011;
DRAM[63458] = 8'b1100100;
DRAM[63459] = 8'b1100100;
DRAM[63460] = 8'b1100101;
DRAM[63461] = 8'b1100110;
DRAM[63462] = 8'b1100111;
DRAM[63463] = 8'b1100111;
DRAM[63464] = 8'b1101001;
DRAM[63465] = 8'b1101000;
DRAM[63466] = 8'b1101000;
DRAM[63467] = 8'b1100111;
DRAM[63468] = 8'b1100111;
DRAM[63469] = 8'b1101000;
DRAM[63470] = 8'b1101000;
DRAM[63471] = 8'b1101001;
DRAM[63472] = 8'b1101000;
DRAM[63473] = 8'b1101010;
DRAM[63474] = 8'b1101101;
DRAM[63475] = 8'b1101111;
DRAM[63476] = 8'b1110000;
DRAM[63477] = 8'b1101111;
DRAM[63478] = 8'b1101110;
DRAM[63479] = 8'b1101101;
DRAM[63480] = 8'b1101100;
DRAM[63481] = 8'b1101100;
DRAM[63482] = 8'b1101011;
DRAM[63483] = 8'b1101010;
DRAM[63484] = 8'b1101001;
DRAM[63485] = 8'b1100111;
DRAM[63486] = 8'b1100111;
DRAM[63487] = 8'b1100110;
DRAM[63488] = 8'b10010011;
DRAM[63489] = 8'b10001101;
DRAM[63490] = 8'b10001101;
DRAM[63491] = 8'b10001111;
DRAM[63492] = 8'b10001101;
DRAM[63493] = 8'b10001110;
DRAM[63494] = 8'b10100000;
DRAM[63495] = 8'b10110111;
DRAM[63496] = 8'b11010011;
DRAM[63497] = 8'b11100101;
DRAM[63498] = 8'b11110011;
DRAM[63499] = 8'b11110010;
DRAM[63500] = 8'b11110010;
DRAM[63501] = 8'b11110111;
DRAM[63502] = 8'b11110101;
DRAM[63503] = 8'b11101110;
DRAM[63504] = 8'b11100101;
DRAM[63505] = 8'b11100111;
DRAM[63506] = 8'b11101001;
DRAM[63507] = 8'b11101100;
DRAM[63508] = 8'b11101100;
DRAM[63509] = 8'b11101000;
DRAM[63510] = 8'b11100001;
DRAM[63511] = 8'b11011100;
DRAM[63512] = 8'b11011011;
DRAM[63513] = 8'b11011000;
DRAM[63514] = 8'b11010100;
DRAM[63515] = 8'b11010001;
DRAM[63516] = 8'b11010000;
DRAM[63517] = 8'b11001110;
DRAM[63518] = 8'b11001100;
DRAM[63519] = 8'b11001010;
DRAM[63520] = 8'b10111110;
DRAM[63521] = 8'b10111101;
DRAM[63522] = 8'b10111010;
DRAM[63523] = 8'b10111011;
DRAM[63524] = 8'b11000011;
DRAM[63525] = 8'b11001010;
DRAM[63526] = 8'b11000110;
DRAM[63527] = 8'b10111110;
DRAM[63528] = 8'b10111010;
DRAM[63529] = 8'b10110011;
DRAM[63530] = 8'b10110001;
DRAM[63531] = 8'b10110100;
DRAM[63532] = 8'b10110101;
DRAM[63533] = 8'b10101111;
DRAM[63534] = 8'b10101110;
DRAM[63535] = 8'b10110000;
DRAM[63536] = 8'b10101011;
DRAM[63537] = 8'b10101001;
DRAM[63538] = 8'b10100101;
DRAM[63539] = 8'b10011111;
DRAM[63540] = 8'b10011001;
DRAM[63541] = 8'b10010011;
DRAM[63542] = 8'b10001110;
DRAM[63543] = 8'b10001100;
DRAM[63544] = 8'b10010100;
DRAM[63545] = 8'b10010001;
DRAM[63546] = 8'b10001111;
DRAM[63547] = 8'b10001111;
DRAM[63548] = 8'b10010011;
DRAM[63549] = 8'b10011000;
DRAM[63550] = 8'b10011100;
DRAM[63551] = 8'b10011110;
DRAM[63552] = 8'b10011011;
DRAM[63553] = 8'b10011101;
DRAM[63554] = 8'b10010011;
DRAM[63555] = 8'b10000010;
DRAM[63556] = 8'b1111111;
DRAM[63557] = 8'b10000110;
DRAM[63558] = 8'b10000000;
DRAM[63559] = 8'b1101111;
DRAM[63560] = 8'b1111100;
DRAM[63561] = 8'b1111110;
DRAM[63562] = 8'b10000001;
DRAM[63563] = 8'b10000010;
DRAM[63564] = 8'b10000001;
DRAM[63565] = 8'b1111110;
DRAM[63566] = 8'b1111010;
DRAM[63567] = 8'b1110111;
DRAM[63568] = 8'b1111111;
DRAM[63569] = 8'b10001000;
DRAM[63570] = 8'b10000111;
DRAM[63571] = 8'b1111100;
DRAM[63572] = 8'b1110111;
DRAM[63573] = 8'b1111100;
DRAM[63574] = 8'b1111111;
DRAM[63575] = 8'b1111101;
DRAM[63576] = 8'b1111000;
DRAM[63577] = 8'b1110001;
DRAM[63578] = 8'b1110110;
DRAM[63579] = 8'b1101111;
DRAM[63580] = 8'b1110101;
DRAM[63581] = 8'b10000010;
DRAM[63582] = 8'b1110100;
DRAM[63583] = 8'b1101111;
DRAM[63584] = 8'b1110101;
DRAM[63585] = 8'b1100111;
DRAM[63586] = 8'b1100101;
DRAM[63587] = 8'b1110100;
DRAM[63588] = 8'b1111100;
DRAM[63589] = 8'b1110111;
DRAM[63590] = 8'b1110110;
DRAM[63591] = 8'b1111101;
DRAM[63592] = 8'b1111110;
DRAM[63593] = 8'b1111011;
DRAM[63594] = 8'b1110100;
DRAM[63595] = 8'b1101111;
DRAM[63596] = 8'b1110011;
DRAM[63597] = 8'b1110111;
DRAM[63598] = 8'b1101111;
DRAM[63599] = 8'b1100010;
DRAM[63600] = 8'b1110011;
DRAM[63601] = 8'b1101001;
DRAM[63602] = 8'b1100010;
DRAM[63603] = 8'b1101001;
DRAM[63604] = 8'b1111001;
DRAM[63605] = 8'b10000001;
DRAM[63606] = 8'b1111011;
DRAM[63607] = 8'b1110000;
DRAM[63608] = 8'b1110100;
DRAM[63609] = 8'b1110001;
DRAM[63610] = 8'b1101101;
DRAM[63611] = 8'b1101100;
DRAM[63612] = 8'b1101011;
DRAM[63613] = 8'b1100110;
DRAM[63614] = 8'b1011111;
DRAM[63615] = 8'b1011001;
DRAM[63616] = 8'b1110101;
DRAM[63617] = 8'b1110100;
DRAM[63618] = 8'b1100000;
DRAM[63619] = 8'b1100010;
DRAM[63620] = 8'b1110111;
DRAM[63621] = 8'b1101100;
DRAM[63622] = 8'b1100001;
DRAM[63623] = 8'b1111010;
DRAM[63624] = 8'b1110000;
DRAM[63625] = 8'b1101111;
DRAM[63626] = 8'b1101111;
DRAM[63627] = 8'b1100111;
DRAM[63628] = 8'b1011100;
DRAM[63629] = 8'b1100101;
DRAM[63630] = 8'b1110010;
DRAM[63631] = 8'b1110000;
DRAM[63632] = 8'b1101110;
DRAM[63633] = 8'b1110000;
DRAM[63634] = 8'b1101110;
DRAM[63635] = 8'b1111000;
DRAM[63636] = 8'b1110010;
DRAM[63637] = 8'b1101100;
DRAM[63638] = 8'b1110110;
DRAM[63639] = 8'b1101000;
DRAM[63640] = 8'b1101110;
DRAM[63641] = 8'b1111010;
DRAM[63642] = 8'b10000000;
DRAM[63643] = 8'b1111000;
DRAM[63644] = 8'b1110011;
DRAM[63645] = 8'b1110110;
DRAM[63646] = 8'b1111001;
DRAM[63647] = 8'b1110110;
DRAM[63648] = 8'b1110010;
DRAM[63649] = 8'b1110111;
DRAM[63650] = 8'b1111101;
DRAM[63651] = 8'b10000000;
DRAM[63652] = 8'b10000000;
DRAM[63653] = 8'b10000001;
DRAM[63654] = 8'b10000011;
DRAM[63655] = 8'b10000110;
DRAM[63656] = 8'b10000011;
DRAM[63657] = 8'b10001001;
DRAM[63658] = 8'b10001100;
DRAM[63659] = 8'b10001100;
DRAM[63660] = 8'b10010000;
DRAM[63661] = 8'b10010110;
DRAM[63662] = 8'b10010100;
DRAM[63663] = 8'b10001101;
DRAM[63664] = 8'b10011011;
DRAM[63665] = 8'b10100000;
DRAM[63666] = 8'b10100010;
DRAM[63667] = 8'b10011110;
DRAM[63668] = 8'b10010111;
DRAM[63669] = 8'b10010101;
DRAM[63670] = 8'b10011000;
DRAM[63671] = 8'b10011110;
DRAM[63672] = 8'b10011110;
DRAM[63673] = 8'b10100001;
DRAM[63674] = 8'b10101001;
DRAM[63675] = 8'b10110100;
DRAM[63676] = 8'b10111110;
DRAM[63677] = 8'b11001001;
DRAM[63678] = 8'b11011011;
DRAM[63679] = 8'b11101011;
DRAM[63680] = 8'b11101011;
DRAM[63681] = 8'b11100000;
DRAM[63682] = 8'b10111100;
DRAM[63683] = 8'b10011100;
DRAM[63684] = 8'b10010110;
DRAM[63685] = 8'b10010101;
DRAM[63686] = 8'b10001101;
DRAM[63687] = 8'b10001001;
DRAM[63688] = 8'b10001000;
DRAM[63689] = 8'b10000001;
DRAM[63690] = 8'b1111100;
DRAM[63691] = 8'b1111011;
DRAM[63692] = 8'b1111000;
DRAM[63693] = 8'b1110010;
DRAM[63694] = 8'b1101111;
DRAM[63695] = 8'b1101111;
DRAM[63696] = 8'b1101011;
DRAM[63697] = 8'b1101001;
DRAM[63698] = 8'b1100110;
DRAM[63699] = 8'b1100011;
DRAM[63700] = 8'b1100000;
DRAM[63701] = 8'b1011101;
DRAM[63702] = 8'b1011100;
DRAM[63703] = 8'b1011011;
DRAM[63704] = 8'b1011101;
DRAM[63705] = 8'b1011101;
DRAM[63706] = 8'b1011101;
DRAM[63707] = 8'b1011110;
DRAM[63708] = 8'b1100000;
DRAM[63709] = 8'b1100010;
DRAM[63710] = 8'b1100100;
DRAM[63711] = 8'b1100101;
DRAM[63712] = 8'b1100001;
DRAM[63713] = 8'b1100010;
DRAM[63714] = 8'b1100011;
DRAM[63715] = 8'b1100100;
DRAM[63716] = 8'b1100101;
DRAM[63717] = 8'b1100110;
DRAM[63718] = 8'b1100101;
DRAM[63719] = 8'b1100101;
DRAM[63720] = 8'b1100110;
DRAM[63721] = 8'b1100110;
DRAM[63722] = 8'b1100110;
DRAM[63723] = 8'b1100111;
DRAM[63724] = 8'b1100111;
DRAM[63725] = 8'b1101000;
DRAM[63726] = 8'b1101000;
DRAM[63727] = 8'b1101000;
DRAM[63728] = 8'b1101010;
DRAM[63729] = 8'b1101011;
DRAM[63730] = 8'b1101100;
DRAM[63731] = 8'b1101101;
DRAM[63732] = 8'b1101101;
DRAM[63733] = 8'b1101101;
DRAM[63734] = 8'b1101101;
DRAM[63735] = 8'b1101100;
DRAM[63736] = 8'b1101100;
DRAM[63737] = 8'b1101100;
DRAM[63738] = 8'b1101011;
DRAM[63739] = 8'b1101010;
DRAM[63740] = 8'b1101000;
DRAM[63741] = 8'b1100111;
DRAM[63742] = 8'b1100110;
DRAM[63743] = 8'b1100110;
DRAM[63744] = 8'b10010010;
DRAM[63745] = 8'b10001101;
DRAM[63746] = 8'b10001011;
DRAM[63747] = 8'b10001101;
DRAM[63748] = 8'b10001100;
DRAM[63749] = 8'b10010000;
DRAM[63750] = 8'b10100011;
DRAM[63751] = 8'b10111011;
DRAM[63752] = 8'b11010101;
DRAM[63753] = 8'b11100110;
DRAM[63754] = 8'b11110001;
DRAM[63755] = 8'b11110000;
DRAM[63756] = 8'b11101111;
DRAM[63757] = 8'b11110011;
DRAM[63758] = 8'b11110001;
DRAM[63759] = 8'b11101010;
DRAM[63760] = 8'b11100100;
DRAM[63761] = 8'b11100101;
DRAM[63762] = 8'b11100111;
DRAM[63763] = 8'b11101010;
DRAM[63764] = 8'b11101010;
DRAM[63765] = 8'b11100110;
DRAM[63766] = 8'b11011111;
DRAM[63767] = 8'b11011001;
DRAM[63768] = 8'b11010011;
DRAM[63769] = 8'b11010001;
DRAM[63770] = 8'b11001101;
DRAM[63771] = 8'b11001011;
DRAM[63772] = 8'b11001001;
DRAM[63773] = 8'b11001000;
DRAM[63774] = 8'b11000101;
DRAM[63775] = 8'b11000011;
DRAM[63776] = 8'b10111010;
DRAM[63777] = 8'b10111010;
DRAM[63778] = 8'b10111000;
DRAM[63779] = 8'b10110111;
DRAM[63780] = 8'b10111100;
DRAM[63781] = 8'b11000010;
DRAM[63782] = 8'b11000001;
DRAM[63783] = 8'b10111100;
DRAM[63784] = 8'b10111010;
DRAM[63785] = 8'b10110010;
DRAM[63786] = 8'b10101100;
DRAM[63787] = 8'b10101011;
DRAM[63788] = 8'b10101001;
DRAM[63789] = 8'b10100101;
DRAM[63790] = 8'b10100100;
DRAM[63791] = 8'b10100110;
DRAM[63792] = 8'b10100110;
DRAM[63793] = 8'b10100100;
DRAM[63794] = 8'b10100010;
DRAM[63795] = 8'b10100000;
DRAM[63796] = 8'b10011101;
DRAM[63797] = 8'b10011011;
DRAM[63798] = 8'b10011010;
DRAM[63799] = 8'b10011001;
DRAM[63800] = 8'b10010100;
DRAM[63801] = 8'b10010000;
DRAM[63802] = 8'b10001100;
DRAM[63803] = 8'b10001110;
DRAM[63804] = 8'b10010100;
DRAM[63805] = 8'b10011010;
DRAM[63806] = 8'b10011100;
DRAM[63807] = 8'b10011100;
DRAM[63808] = 8'b10010001;
DRAM[63809] = 8'b10010101;
DRAM[63810] = 8'b10010010;
DRAM[63811] = 8'b10001001;
DRAM[63812] = 8'b10000111;
DRAM[63813] = 8'b10001000;
DRAM[63814] = 8'b10000000;
DRAM[63815] = 8'b1110011;
DRAM[63816] = 8'b10000001;
DRAM[63817] = 8'b1111110;
DRAM[63818] = 8'b1111001;
DRAM[63819] = 8'b1110101;
DRAM[63820] = 8'b1110011;
DRAM[63821] = 8'b1110101;
DRAM[63822] = 8'b1111000;
DRAM[63823] = 8'b1111011;
DRAM[63824] = 8'b1101000;
DRAM[63825] = 8'b1101100;
DRAM[63826] = 8'b1110000;
DRAM[63827] = 8'b1110110;
DRAM[63828] = 8'b1111110;
DRAM[63829] = 8'b10000010;
DRAM[63830] = 8'b1111101;
DRAM[63831] = 8'b1110100;
DRAM[63832] = 8'b1111001;
DRAM[63833] = 8'b1110011;
DRAM[63834] = 8'b1110111;
DRAM[63835] = 8'b1101110;
DRAM[63836] = 8'b1110010;
DRAM[63837] = 8'b1111110;
DRAM[63838] = 8'b1110010;
DRAM[63839] = 8'b1110001;
DRAM[63840] = 8'b1101111;
DRAM[63841] = 8'b1100101;
DRAM[63842] = 8'b1101000;
DRAM[63843] = 8'b1110110;
DRAM[63844] = 8'b1111011;
DRAM[63845] = 8'b1110010;
DRAM[63846] = 8'b1101111;
DRAM[63847] = 8'b1110101;
DRAM[63848] = 8'b1111001;
DRAM[63849] = 8'b1111010;
DRAM[63850] = 8'b1111101;
DRAM[63851] = 8'b1111110;
DRAM[63852] = 8'b1110101;
DRAM[63853] = 8'b1101010;
DRAM[63854] = 8'b1101011;
DRAM[63855] = 8'b1110100;
DRAM[63856] = 8'b1110111;
DRAM[63857] = 8'b1110000;
DRAM[63858] = 8'b1101001;
DRAM[63859] = 8'b1101000;
DRAM[63860] = 8'b1101100;
DRAM[63861] = 8'b1110000;
DRAM[63862] = 8'b1101111;
DRAM[63863] = 8'b1101100;
DRAM[63864] = 8'b1110101;
DRAM[63865] = 8'b1110101;
DRAM[63866] = 8'b1110100;
DRAM[63867] = 8'b1110101;
DRAM[63868] = 8'b1110101;
DRAM[63869] = 8'b1110100;
DRAM[63870] = 8'b1110001;
DRAM[63871] = 8'b1101111;
DRAM[63872] = 8'b1100101;
DRAM[63873] = 8'b1101101;
DRAM[63874] = 8'b1100000;
DRAM[63875] = 8'b1011010;
DRAM[63876] = 8'b1101010;
DRAM[63877] = 8'b1101110;
DRAM[63878] = 8'b1101000;
DRAM[63879] = 8'b1101110;
DRAM[63880] = 8'b1101110;
DRAM[63881] = 8'b1101110;
DRAM[63882] = 8'b1110001;
DRAM[63883] = 8'b1101011;
DRAM[63884] = 8'b1100000;
DRAM[63885] = 8'b1100111;
DRAM[63886] = 8'b1110011;
DRAM[63887] = 8'b1110001;
DRAM[63888] = 8'b1101100;
DRAM[63889] = 8'b1101110;
DRAM[63890] = 8'b1101100;
DRAM[63891] = 8'b1110111;
DRAM[63892] = 8'b1110010;
DRAM[63893] = 8'b1101110;
DRAM[63894] = 8'b1111001;
DRAM[63895] = 8'b1101011;
DRAM[63896] = 8'b1100111;
DRAM[63897] = 8'b1110010;
DRAM[63898] = 8'b1111011;
DRAM[63899] = 8'b1111011;
DRAM[63900] = 8'b1111000;
DRAM[63901] = 8'b1111000;
DRAM[63902] = 8'b1111000;
DRAM[63903] = 8'b1110111;
DRAM[63904] = 8'b1110010;
DRAM[63905] = 8'b1110101;
DRAM[63906] = 8'b1111010;
DRAM[63907] = 8'b1111101;
DRAM[63908] = 8'b1111111;
DRAM[63909] = 8'b10000001;
DRAM[63910] = 8'b10000011;
DRAM[63911] = 8'b10000100;
DRAM[63912] = 8'b10000001;
DRAM[63913] = 8'b10000110;
DRAM[63914] = 8'b10001001;
DRAM[63915] = 8'b10001011;
DRAM[63916] = 8'b10001111;
DRAM[63917] = 8'b10010101;
DRAM[63918] = 8'b10010100;
DRAM[63919] = 8'b10001110;
DRAM[63920] = 8'b10010000;
DRAM[63921] = 8'b10010100;
DRAM[63922] = 8'b10011000;
DRAM[63923] = 8'b10010110;
DRAM[63924] = 8'b10010010;
DRAM[63925] = 8'b10010001;
DRAM[63926] = 8'b10010111;
DRAM[63927] = 8'b10011110;
DRAM[63928] = 8'b10100111;
DRAM[63929] = 8'b10101010;
DRAM[63930] = 8'b10110001;
DRAM[63931] = 8'b10111011;
DRAM[63932] = 8'b11000011;
DRAM[63933] = 8'b11001101;
DRAM[63934] = 8'b11011100;
DRAM[63935] = 8'b11101010;
DRAM[63936] = 8'b11101101;
DRAM[63937] = 8'b11100111;
DRAM[63938] = 8'b11001000;
DRAM[63939] = 8'b10100100;
DRAM[63940] = 8'b10010110;
DRAM[63941] = 8'b10010000;
DRAM[63942] = 8'b10001010;
DRAM[63943] = 8'b10001010;
DRAM[63944] = 8'b10000110;
DRAM[63945] = 8'b10000000;
DRAM[63946] = 8'b1111011;
DRAM[63947] = 8'b1111010;
DRAM[63948] = 8'b1110111;
DRAM[63949] = 8'b1110000;
DRAM[63950] = 8'b1101100;
DRAM[63951] = 8'b1101011;
DRAM[63952] = 8'b1101001;
DRAM[63953] = 8'b1101000;
DRAM[63954] = 8'b1100101;
DRAM[63955] = 8'b1100010;
DRAM[63956] = 8'b1011111;
DRAM[63957] = 8'b1011101;
DRAM[63958] = 8'b1011100;
DRAM[63959] = 8'b1011011;
DRAM[63960] = 8'b1011011;
DRAM[63961] = 8'b1011011;
DRAM[63962] = 8'b1011100;
DRAM[63963] = 8'b1011101;
DRAM[63964] = 8'b1011111;
DRAM[63965] = 8'b1100001;
DRAM[63966] = 8'b1100010;
DRAM[63967] = 8'b1100100;
DRAM[63968] = 8'b1100001;
DRAM[63969] = 8'b1100010;
DRAM[63970] = 8'b1100011;
DRAM[63971] = 8'b1100100;
DRAM[63972] = 8'b1100101;
DRAM[63973] = 8'b1100110;
DRAM[63974] = 8'b1100101;
DRAM[63975] = 8'b1100101;
DRAM[63976] = 8'b1100110;
DRAM[63977] = 8'b1100110;
DRAM[63978] = 8'b1100110;
DRAM[63979] = 8'b1100111;
DRAM[63980] = 8'b1100111;
DRAM[63981] = 8'b1101000;
DRAM[63982] = 8'b1101000;
DRAM[63983] = 8'b1101000;
DRAM[63984] = 8'b1101010;
DRAM[63985] = 8'b1101011;
DRAM[63986] = 8'b1101100;
DRAM[63987] = 8'b1101100;
DRAM[63988] = 8'b1101101;
DRAM[63989] = 8'b1101101;
DRAM[63990] = 8'b1101100;
DRAM[63991] = 8'b1101100;
DRAM[63992] = 8'b1101100;
DRAM[63993] = 8'b1101100;
DRAM[63994] = 8'b1101011;
DRAM[63995] = 8'b1101010;
DRAM[63996] = 8'b1101000;
DRAM[63997] = 8'b1100111;
DRAM[63998] = 8'b1100110;
DRAM[63999] = 8'b1100110;
DRAM[64000] = 8'b10010101;
DRAM[64001] = 8'b10001111;
DRAM[64002] = 8'b10001100;
DRAM[64003] = 8'b10001101;
DRAM[64004] = 8'b10001110;
DRAM[64005] = 8'b10010110;
DRAM[64006] = 8'b10101100;
DRAM[64007] = 8'b11000100;
DRAM[64008] = 8'b11011010;
DRAM[64009] = 8'b11100111;
DRAM[64010] = 8'b11101111;
DRAM[64011] = 8'b11101110;
DRAM[64012] = 8'b11101100;
DRAM[64013] = 8'b11101101;
DRAM[64014] = 8'b11101011;
DRAM[64015] = 8'b11100100;
DRAM[64016] = 8'b11100010;
DRAM[64017] = 8'b11100011;
DRAM[64018] = 8'b11100101;
DRAM[64019] = 8'b11101000;
DRAM[64020] = 8'b11100111;
DRAM[64021] = 8'b11100011;
DRAM[64022] = 8'b11011100;
DRAM[64023] = 8'b11010110;
DRAM[64024] = 8'b11010100;
DRAM[64025] = 8'b11010001;
DRAM[64026] = 8'b11001110;
DRAM[64027] = 8'b11001100;
DRAM[64028] = 8'b11001011;
DRAM[64029] = 8'b11001001;
DRAM[64030] = 8'b11000110;
DRAM[64031] = 8'b11000011;
DRAM[64032] = 8'b11000110;
DRAM[64033] = 8'b11000110;
DRAM[64034] = 8'b11000011;
DRAM[64035] = 8'b10111110;
DRAM[64036] = 8'b10111101;
DRAM[64037] = 8'b10111111;
DRAM[64038] = 8'b10111100;
DRAM[64039] = 8'b10110110;
DRAM[64040] = 8'b10110111;
DRAM[64041] = 8'b10101111;
DRAM[64042] = 8'b10100111;
DRAM[64043] = 8'b10100011;
DRAM[64044] = 8'b10100001;
DRAM[64045] = 8'b10011110;
DRAM[64046] = 8'b10011110;
DRAM[64047] = 8'b10100001;
DRAM[64048] = 8'b10100110;
DRAM[64049] = 8'b10100110;
DRAM[64050] = 8'b10100101;
DRAM[64051] = 8'b10100101;
DRAM[64052] = 8'b10100100;
DRAM[64053] = 8'b10100100;
DRAM[64054] = 8'b10100100;
DRAM[64055] = 8'b10100100;
DRAM[64056] = 8'b10011100;
DRAM[64057] = 8'b10010111;
DRAM[64058] = 8'b10010010;
DRAM[64059] = 8'b10010010;
DRAM[64060] = 8'b10010101;
DRAM[64061] = 8'b10010110;
DRAM[64062] = 8'b10010011;
DRAM[64063] = 8'b10010000;
DRAM[64064] = 8'b10001110;
DRAM[64065] = 8'b10001101;
DRAM[64066] = 8'b10001010;
DRAM[64067] = 8'b10000110;
DRAM[64068] = 8'b10000000;
DRAM[64069] = 8'b1111010;
DRAM[64070] = 8'b1110101;
DRAM[64071] = 8'b1110001;
DRAM[64072] = 8'b1101111;
DRAM[64073] = 8'b1110000;
DRAM[64074] = 8'b1110001;
DRAM[64075] = 8'b1110010;
DRAM[64076] = 8'b1110001;
DRAM[64077] = 8'b1101111;
DRAM[64078] = 8'b1101101;
DRAM[64079] = 8'b1101011;
DRAM[64080] = 8'b1101011;
DRAM[64081] = 8'b1101000;
DRAM[64082] = 8'b1101010;
DRAM[64083] = 8'b1110010;
DRAM[64084] = 8'b1111000;
DRAM[64085] = 8'b1111010;
DRAM[64086] = 8'b1111010;
DRAM[64087] = 8'b1111011;
DRAM[64088] = 8'b1111100;
DRAM[64089] = 8'b1110100;
DRAM[64090] = 8'b1111000;
DRAM[64091] = 8'b1101101;
DRAM[64092] = 8'b1101101;
DRAM[64093] = 8'b1110111;
DRAM[64094] = 8'b1101111;
DRAM[64095] = 8'b1110010;
DRAM[64096] = 8'b1101010;
DRAM[64097] = 8'b1100100;
DRAM[64098] = 8'b1101001;
DRAM[64099] = 8'b1111000;
DRAM[64100] = 8'b1111011;
DRAM[64101] = 8'b1110000;
DRAM[64102] = 8'b1101001;
DRAM[64103] = 8'b1101100;
DRAM[64104] = 8'b1110110;
DRAM[64105] = 8'b1110000;
DRAM[64106] = 8'b1110110;
DRAM[64107] = 8'b1111111;
DRAM[64108] = 8'b1110110;
DRAM[64109] = 8'b1100100;
DRAM[64110] = 8'b1100101;
DRAM[64111] = 8'b1110101;
DRAM[64112] = 8'b1101111;
DRAM[64113] = 8'b1101111;
DRAM[64114] = 8'b1101101;
DRAM[64115] = 8'b1101001;
DRAM[64116] = 8'b1100111;
DRAM[64117] = 8'b1101011;
DRAM[64118] = 8'b1110011;
DRAM[64119] = 8'b1111011;
DRAM[64120] = 8'b1101010;
DRAM[64121] = 8'b1101011;
DRAM[64122] = 8'b1101011;
DRAM[64123] = 8'b1101010;
DRAM[64124] = 8'b1101001;
DRAM[64125] = 8'b1101001;
DRAM[64126] = 8'b1101010;
DRAM[64127] = 8'b1101011;
DRAM[64128] = 8'b1100101;
DRAM[64129] = 8'b1101111;
DRAM[64130] = 8'b1101010;
DRAM[64131] = 8'b1011100;
DRAM[64132] = 8'b1100010;
DRAM[64133] = 8'b1110101;
DRAM[64134] = 8'b1110110;
DRAM[64135] = 8'b1101001;
DRAM[64136] = 8'b1101010;
DRAM[64137] = 8'b1101100;
DRAM[64138] = 8'b1110011;
DRAM[64139] = 8'b1110000;
DRAM[64140] = 8'b1100101;
DRAM[64141] = 8'b1101001;
DRAM[64142] = 8'b1110100;
DRAM[64143] = 8'b1110011;
DRAM[64144] = 8'b1101011;
DRAM[64145] = 8'b1101100;
DRAM[64146] = 8'b1101001;
DRAM[64147] = 8'b1110101;
DRAM[64148] = 8'b1110011;
DRAM[64149] = 8'b1110000;
DRAM[64150] = 8'b1111100;
DRAM[64151] = 8'b1101110;
DRAM[64152] = 8'b1100011;
DRAM[64153] = 8'b1101001;
DRAM[64154] = 8'b1110100;
DRAM[64155] = 8'b1111110;
DRAM[64156] = 8'b1111110;
DRAM[64157] = 8'b1111001;
DRAM[64158] = 8'b1110111;
DRAM[64159] = 8'b1111001;
DRAM[64160] = 8'b1110011;
DRAM[64161] = 8'b1110011;
DRAM[64162] = 8'b1110101;
DRAM[64163] = 8'b1111001;
DRAM[64164] = 8'b1111101;
DRAM[64165] = 8'b10000001;
DRAM[64166] = 8'b10000010;
DRAM[64167] = 8'b10000010;
DRAM[64168] = 8'b10000011;
DRAM[64169] = 8'b10000111;
DRAM[64170] = 8'b10001001;
DRAM[64171] = 8'b10001011;
DRAM[64172] = 8'b10001111;
DRAM[64173] = 8'b10010100;
DRAM[64174] = 8'b10010100;
DRAM[64175] = 8'b10010000;
DRAM[64176] = 8'b10001000;
DRAM[64177] = 8'b10001101;
DRAM[64178] = 8'b10010001;
DRAM[64179] = 8'b10010010;
DRAM[64180] = 8'b10010001;
DRAM[64181] = 8'b10010100;
DRAM[64182] = 8'b10011100;
DRAM[64183] = 8'b10100100;
DRAM[64184] = 8'b10101100;
DRAM[64185] = 8'b10101110;
DRAM[64186] = 8'b10110101;
DRAM[64187] = 8'b10111110;
DRAM[64188] = 8'b11000101;
DRAM[64189] = 8'b11001100;
DRAM[64190] = 8'b11010111;
DRAM[64191] = 8'b11100011;
DRAM[64192] = 8'b11101101;
DRAM[64193] = 8'b11101011;
DRAM[64194] = 8'b11001101;
DRAM[64195] = 8'b10100100;
DRAM[64196] = 8'b10001111;
DRAM[64197] = 8'b10000110;
DRAM[64198] = 8'b10000100;
DRAM[64199] = 8'b10001010;
DRAM[64200] = 8'b10000000;
DRAM[64201] = 8'b1111011;
DRAM[64202] = 8'b1111000;
DRAM[64203] = 8'b1111000;
DRAM[64204] = 8'b1110110;
DRAM[64205] = 8'b1101111;
DRAM[64206] = 8'b1101011;
DRAM[64207] = 8'b1101010;
DRAM[64208] = 8'b1100111;
DRAM[64209] = 8'b1100101;
DRAM[64210] = 8'b1100011;
DRAM[64211] = 8'b1100001;
DRAM[64212] = 8'b1011110;
DRAM[64213] = 8'b1011101;
DRAM[64214] = 8'b1011100;
DRAM[64215] = 8'b1011100;
DRAM[64216] = 8'b1011010;
DRAM[64217] = 8'b1011010;
DRAM[64218] = 8'b1011010;
DRAM[64219] = 8'b1011011;
DRAM[64220] = 8'b1011101;
DRAM[64221] = 8'b1011111;
DRAM[64222] = 8'b1100001;
DRAM[64223] = 8'b1100010;
DRAM[64224] = 8'b1100001;
DRAM[64225] = 8'b1100010;
DRAM[64226] = 8'b1100011;
DRAM[64227] = 8'b1100100;
DRAM[64228] = 8'b1100101;
DRAM[64229] = 8'b1100110;
DRAM[64230] = 8'b1100101;
DRAM[64231] = 8'b1100101;
DRAM[64232] = 8'b1100110;
DRAM[64233] = 8'b1100110;
DRAM[64234] = 8'b1100110;
DRAM[64235] = 8'b1100111;
DRAM[64236] = 8'b1100111;
DRAM[64237] = 8'b1101000;
DRAM[64238] = 8'b1101000;
DRAM[64239] = 8'b1101000;
DRAM[64240] = 8'b1101010;
DRAM[64241] = 8'b1101010;
DRAM[64242] = 8'b1101011;
DRAM[64243] = 8'b1101100;
DRAM[64244] = 8'b1101101;
DRAM[64245] = 8'b1101101;
DRAM[64246] = 8'b1101100;
DRAM[64247] = 8'b1101100;
DRAM[64248] = 8'b1101100;
DRAM[64249] = 8'b1101100;
DRAM[64250] = 8'b1101011;
DRAM[64251] = 8'b1101010;
DRAM[64252] = 8'b1101000;
DRAM[64253] = 8'b1100111;
DRAM[64254] = 8'b1100110;
DRAM[64255] = 8'b1100110;
DRAM[64256] = 8'b10010111;
DRAM[64257] = 8'b10010001;
DRAM[64258] = 8'b10001110;
DRAM[64259] = 8'b10001111;
DRAM[64260] = 8'b10010011;
DRAM[64261] = 8'b10100000;
DRAM[64262] = 8'b10111001;
DRAM[64263] = 8'b11001111;
DRAM[64264] = 8'b11100001;
DRAM[64265] = 8'b11101001;
DRAM[64266] = 8'b11101110;
DRAM[64267] = 8'b11101100;
DRAM[64268] = 8'b11101001;
DRAM[64269] = 8'b11101001;
DRAM[64270] = 8'b11100101;
DRAM[64271] = 8'b11100000;
DRAM[64272] = 8'b11100001;
DRAM[64273] = 8'b11100010;
DRAM[64274] = 8'b11100100;
DRAM[64275] = 8'b11100110;
DRAM[64276] = 8'b11100110;
DRAM[64277] = 8'b11100001;
DRAM[64278] = 8'b11011010;
DRAM[64279] = 8'b11010101;
DRAM[64280] = 8'b11010110;
DRAM[64281] = 8'b11010100;
DRAM[64282] = 8'b11010001;
DRAM[64283] = 8'b11010000;
DRAM[64284] = 8'b11001110;
DRAM[64285] = 8'b11001100;
DRAM[64286] = 8'b11001000;
DRAM[64287] = 8'b11000101;
DRAM[64288] = 8'b11001001;
DRAM[64289] = 8'b11001000;
DRAM[64290] = 8'b11000110;
DRAM[64291] = 8'b11000011;
DRAM[64292] = 8'b11000101;
DRAM[64293] = 8'b11000101;
DRAM[64294] = 8'b10111101;
DRAM[64295] = 8'b10110011;
DRAM[64296] = 8'b10110010;
DRAM[64297] = 8'b10101100;
DRAM[64298] = 8'b10100110;
DRAM[64299] = 8'b10100011;
DRAM[64300] = 8'b10100010;
DRAM[64301] = 8'b10100001;
DRAM[64302] = 8'b10100001;
DRAM[64303] = 8'b10100010;
DRAM[64304] = 8'b10100100;
DRAM[64305] = 8'b10100101;
DRAM[64306] = 8'b10100110;
DRAM[64307] = 8'b10100101;
DRAM[64308] = 8'b10100011;
DRAM[64309] = 8'b10100000;
DRAM[64310] = 8'b10011101;
DRAM[64311] = 8'b10011011;
DRAM[64312] = 8'b10011000;
DRAM[64313] = 8'b10011000;
DRAM[64314] = 8'b10011001;
DRAM[64315] = 8'b10011001;
DRAM[64316] = 8'b10010111;
DRAM[64317] = 8'b10010100;
DRAM[64318] = 8'b10010000;
DRAM[64319] = 8'b10001101;
DRAM[64320] = 8'b10001111;
DRAM[64321] = 8'b10000110;
DRAM[64322] = 8'b1111111;
DRAM[64323] = 8'b1111101;
DRAM[64324] = 8'b1111000;
DRAM[64325] = 8'b1110001;
DRAM[64326] = 8'b1110100;
DRAM[64327] = 8'b1111101;
DRAM[64328] = 8'b1101010;
DRAM[64329] = 8'b1101100;
DRAM[64330] = 8'b1101111;
DRAM[64331] = 8'b1110000;
DRAM[64332] = 8'b1110000;
DRAM[64333] = 8'b1101101;
DRAM[64334] = 8'b1101001;
DRAM[64335] = 8'b1100110;
DRAM[64336] = 8'b1101010;
DRAM[64337] = 8'b1101001;
DRAM[64338] = 8'b1101111;
DRAM[64339] = 8'b1110101;
DRAM[64340] = 8'b1110010;
DRAM[64341] = 8'b1101101;
DRAM[64342] = 8'b1110011;
DRAM[64343] = 8'b10000001;
DRAM[64344] = 8'b1111101;
DRAM[64345] = 8'b1110100;
DRAM[64346] = 8'b1110111;
DRAM[64347] = 8'b1101100;
DRAM[64348] = 8'b1101010;
DRAM[64349] = 8'b1110010;
DRAM[64350] = 8'b1101100;
DRAM[64351] = 8'b1110010;
DRAM[64352] = 8'b1101100;
DRAM[64353] = 8'b1100101;
DRAM[64354] = 8'b1100111;
DRAM[64355] = 8'b1110101;
DRAM[64356] = 8'b1111100;
DRAM[64357] = 8'b1110100;
DRAM[64358] = 8'b1101011;
DRAM[64359] = 8'b1101001;
DRAM[64360] = 8'b1111001;
DRAM[64361] = 8'b1101011;
DRAM[64362] = 8'b1100111;
DRAM[64363] = 8'b1110011;
DRAM[64364] = 8'b1111001;
DRAM[64365] = 8'b1110001;
DRAM[64366] = 8'b1101001;
DRAM[64367] = 8'b1100111;
DRAM[64368] = 8'b1101000;
DRAM[64369] = 8'b1101010;
DRAM[64370] = 8'b1101011;
DRAM[64371] = 8'b1101000;
DRAM[64372] = 8'b1100101;
DRAM[64373] = 8'b1101001;
DRAM[64374] = 8'b1110100;
DRAM[64375] = 8'b1111101;
DRAM[64376] = 8'b10000100;
DRAM[64377] = 8'b10000101;
DRAM[64378] = 8'b10000100;
DRAM[64379] = 8'b1111111;
DRAM[64380] = 8'b1111010;
DRAM[64381] = 8'b1111000;
DRAM[64382] = 8'b1111011;
DRAM[64383] = 8'b1111110;
DRAM[64384] = 8'b1110011;
DRAM[64385] = 8'b1110101;
DRAM[64386] = 8'b1110010;
DRAM[64387] = 8'b1100100;
DRAM[64388] = 8'b1100001;
DRAM[64389] = 8'b1110100;
DRAM[64390] = 8'b1111011;
DRAM[64391] = 8'b1101100;
DRAM[64392] = 8'b1100101;
DRAM[64393] = 8'b1100111;
DRAM[64394] = 8'b1110010;
DRAM[64395] = 8'b1110011;
DRAM[64396] = 8'b1101001;
DRAM[64397] = 8'b1101011;
DRAM[64398] = 8'b1110011;
DRAM[64399] = 8'b1110010;
DRAM[64400] = 8'b1101110;
DRAM[64401] = 8'b1101101;
DRAM[64402] = 8'b1101001;
DRAM[64403] = 8'b1110101;
DRAM[64404] = 8'b1110011;
DRAM[64405] = 8'b1110001;
DRAM[64406] = 8'b1111100;
DRAM[64407] = 8'b1101110;
DRAM[64408] = 8'b1100110;
DRAM[64409] = 8'b1100110;
DRAM[64410] = 8'b1110000;
DRAM[64411] = 8'b1111110;
DRAM[64412] = 8'b10000000;
DRAM[64413] = 8'b1111001;
DRAM[64414] = 8'b1110110;
DRAM[64415] = 8'b1111010;
DRAM[64416] = 8'b1110110;
DRAM[64417] = 8'b1110011;
DRAM[64418] = 8'b1110010;
DRAM[64419] = 8'b1110101;
DRAM[64420] = 8'b1111011;
DRAM[64421] = 8'b10000000;
DRAM[64422] = 8'b10000001;
DRAM[64423] = 8'b10000001;
DRAM[64424] = 8'b10000010;
DRAM[64425] = 8'b10000011;
DRAM[64426] = 8'b10000100;
DRAM[64427] = 8'b10000110;
DRAM[64428] = 8'b10001001;
DRAM[64429] = 8'b10001100;
DRAM[64430] = 8'b10001100;
DRAM[64431] = 8'b10001010;
DRAM[64432] = 8'b10000101;
DRAM[64433] = 8'b10001000;
DRAM[64434] = 8'b10001101;
DRAM[64435] = 8'b10001111;
DRAM[64436] = 8'b10010001;
DRAM[64437] = 8'b10010110;
DRAM[64438] = 8'b10011111;
DRAM[64439] = 8'b10100110;
DRAM[64440] = 8'b10101110;
DRAM[64441] = 8'b10110000;
DRAM[64442] = 8'b10110111;
DRAM[64443] = 8'b11000010;
DRAM[64444] = 8'b11001001;
DRAM[64445] = 8'b11001110;
DRAM[64446] = 8'b11010111;
DRAM[64447] = 8'b11100000;
DRAM[64448] = 8'b11101011;
DRAM[64449] = 8'b11101001;
DRAM[64450] = 8'b11001100;
DRAM[64451] = 8'b10100011;
DRAM[64452] = 8'b10001101;
DRAM[64453] = 8'b10000011;
DRAM[64454] = 8'b10000001;
DRAM[64455] = 8'b10000110;
DRAM[64456] = 8'b1111100;
DRAM[64457] = 8'b1110111;
DRAM[64458] = 8'b1110101;
DRAM[64459] = 8'b1110111;
DRAM[64460] = 8'b1110110;
DRAM[64461] = 8'b1110000;
DRAM[64462] = 8'b1101100;
DRAM[64463] = 8'b1101011;
DRAM[64464] = 8'b1100100;
DRAM[64465] = 8'b1100011;
DRAM[64466] = 8'b1100001;
DRAM[64467] = 8'b1011111;
DRAM[64468] = 8'b1011101;
DRAM[64469] = 8'b1011100;
DRAM[64470] = 8'b1011011;
DRAM[64471] = 8'b1011011;
DRAM[64472] = 8'b1011001;
DRAM[64473] = 8'b1011010;
DRAM[64474] = 8'b1011010;
DRAM[64475] = 8'b1011011;
DRAM[64476] = 8'b1011101;
DRAM[64477] = 8'b1011111;
DRAM[64478] = 8'b1100001;
DRAM[64479] = 8'b1100010;
DRAM[64480] = 8'b1100001;
DRAM[64481] = 8'b1100010;
DRAM[64482] = 8'b1100011;
DRAM[64483] = 8'b1100100;
DRAM[64484] = 8'b1100101;
DRAM[64485] = 8'b1100110;
DRAM[64486] = 8'b1100101;
DRAM[64487] = 8'b1100101;
DRAM[64488] = 8'b1100110;
DRAM[64489] = 8'b1100110;
DRAM[64490] = 8'b1100110;
DRAM[64491] = 8'b1100111;
DRAM[64492] = 8'b1100111;
DRAM[64493] = 8'b1101000;
DRAM[64494] = 8'b1101000;
DRAM[64495] = 8'b1101000;
DRAM[64496] = 8'b1101001;
DRAM[64497] = 8'b1101010;
DRAM[64498] = 8'b1101011;
DRAM[64499] = 8'b1101100;
DRAM[64500] = 8'b1101100;
DRAM[64501] = 8'b1101100;
DRAM[64502] = 8'b1101100;
DRAM[64503] = 8'b1101011;
DRAM[64504] = 8'b1101100;
DRAM[64505] = 8'b1101100;
DRAM[64506] = 8'b1101011;
DRAM[64507] = 8'b1101010;
DRAM[64508] = 8'b1101000;
DRAM[64509] = 8'b1100111;
DRAM[64510] = 8'b1100110;
DRAM[64511] = 8'b1100110;
DRAM[64512] = 8'b10010100;
DRAM[64513] = 8'b10010001;
DRAM[64514] = 8'b10001111;
DRAM[64515] = 8'b10010001;
DRAM[64516] = 8'b10011001;
DRAM[64517] = 8'b10101001;
DRAM[64518] = 8'b11000010;
DRAM[64519] = 8'b11010110;
DRAM[64520] = 8'b11100110;
DRAM[64521] = 8'b11101010;
DRAM[64522] = 8'b11101101;
DRAM[64523] = 8'b11101010;
DRAM[64524] = 8'b11100111;
DRAM[64525] = 8'b11100110;
DRAM[64526] = 8'b11100010;
DRAM[64527] = 8'b11011111;
DRAM[64528] = 8'b11100001;
DRAM[64529] = 8'b11100010;
DRAM[64530] = 8'b11100100;
DRAM[64531] = 8'b11100110;
DRAM[64532] = 8'b11100101;
DRAM[64533] = 8'b11100000;
DRAM[64534] = 8'b11011001;
DRAM[64535] = 8'b11010011;
DRAM[64536] = 8'b11010001;
DRAM[64537] = 8'b11010000;
DRAM[64538] = 8'b11001101;
DRAM[64539] = 8'b11001100;
DRAM[64540] = 8'b11001011;
DRAM[64541] = 8'b11001000;
DRAM[64542] = 8'b11000100;
DRAM[64543] = 8'b11000001;
DRAM[64544] = 8'b10111010;
DRAM[64545] = 8'b10111010;
DRAM[64546] = 8'b10111010;
DRAM[64547] = 8'b10111110;
DRAM[64548] = 8'b11000110;
DRAM[64549] = 8'b11001000;
DRAM[64550] = 8'b10111100;
DRAM[64551] = 8'b10101110;
DRAM[64552] = 8'b10101110;
DRAM[64553] = 8'b10101011;
DRAM[64554] = 8'b10100111;
DRAM[64555] = 8'b10100100;
DRAM[64556] = 8'b10100011;
DRAM[64557] = 8'b10100010;
DRAM[64558] = 8'b10100000;
DRAM[64559] = 8'b10011101;
DRAM[64560] = 8'b10011010;
DRAM[64561] = 8'b10011100;
DRAM[64562] = 8'b10011101;
DRAM[64563] = 8'b10011101;
DRAM[64564] = 8'b10011010;
DRAM[64565] = 8'b10010101;
DRAM[64566] = 8'b10001111;
DRAM[64567] = 8'b10001011;
DRAM[64568] = 8'b10001100;
DRAM[64569] = 8'b10010011;
DRAM[64570] = 8'b10011011;
DRAM[64571] = 8'b10011101;
DRAM[64572] = 8'b10011001;
DRAM[64573] = 8'b10010101;
DRAM[64574] = 8'b10010011;
DRAM[64575] = 8'b10010011;
DRAM[64576] = 8'b10001101;
DRAM[64577] = 8'b10000011;
DRAM[64578] = 8'b10000000;
DRAM[64579] = 8'b10000011;
DRAM[64580] = 8'b10000001;
DRAM[64581] = 8'b1111100;
DRAM[64582] = 8'b10000010;
DRAM[64583] = 8'b10001110;
DRAM[64584] = 8'b10000000;
DRAM[64585] = 8'b1111010;
DRAM[64586] = 8'b1110000;
DRAM[64587] = 8'b1101000;
DRAM[64588] = 8'b1100101;
DRAM[64589] = 8'b1100111;
DRAM[64590] = 8'b1101100;
DRAM[64591] = 8'b1110000;
DRAM[64592] = 8'b1011100;
DRAM[64593] = 8'b1011011;
DRAM[64594] = 8'b1100001;
DRAM[64595] = 8'b1101011;
DRAM[64596] = 8'b1101101;
DRAM[64597] = 8'b1101000;
DRAM[64598] = 8'b1101010;
DRAM[64599] = 8'b1110011;
DRAM[64600] = 8'b1111101;
DRAM[64601] = 8'b1110010;
DRAM[64602] = 8'b1110110;
DRAM[64603] = 8'b1101100;
DRAM[64604] = 8'b1101010;
DRAM[64605] = 8'b1101111;
DRAM[64606] = 8'b1101000;
DRAM[64607] = 8'b1110000;
DRAM[64608] = 8'b1110011;
DRAM[64609] = 8'b1100111;
DRAM[64610] = 8'b1100100;
DRAM[64611] = 8'b1110000;
DRAM[64612] = 8'b1111011;
DRAM[64613] = 8'b1111010;
DRAM[64614] = 8'b1110001;
DRAM[64615] = 8'b1101100;
DRAM[64616] = 8'b1111001;
DRAM[64617] = 8'b1110001;
DRAM[64618] = 8'b1101001;
DRAM[64619] = 8'b1101100;
DRAM[64620] = 8'b1111000;
DRAM[64621] = 8'b1111101;
DRAM[64622] = 8'b1110010;
DRAM[64623] = 8'b1100010;
DRAM[64624] = 8'b1101011;
DRAM[64625] = 8'b1101010;
DRAM[64626] = 8'b1100111;
DRAM[64627] = 8'b1100100;
DRAM[64628] = 8'b1100010;
DRAM[64629] = 8'b1100001;
DRAM[64630] = 8'b1100011;
DRAM[64631] = 8'b1100100;
DRAM[64632] = 8'b1101101;
DRAM[64633] = 8'b1101101;
DRAM[64634] = 8'b1101101;
DRAM[64635] = 8'b1101001;
DRAM[64636] = 8'b1100101;
DRAM[64637] = 8'b1100100;
DRAM[64638] = 8'b1101000;
DRAM[64639] = 8'b1101101;
DRAM[64640] = 8'b1111100;
DRAM[64641] = 8'b1110000;
DRAM[64642] = 8'b1101010;
DRAM[64643] = 8'b1100110;
DRAM[64644] = 8'b1100001;
DRAM[64645] = 8'b1101001;
DRAM[64646] = 8'b1110011;
DRAM[64647] = 8'b1110010;
DRAM[64648] = 8'b1100011;
DRAM[64649] = 8'b1100011;
DRAM[64650] = 8'b1101111;
DRAM[64651] = 8'b1110100;
DRAM[64652] = 8'b1101101;
DRAM[64653] = 8'b1101101;
DRAM[64654] = 8'b1110010;
DRAM[64655] = 8'b1101111;
DRAM[64656] = 8'b1110001;
DRAM[64657] = 8'b1110000;
DRAM[64658] = 8'b1101011;
DRAM[64659] = 8'b1110110;
DRAM[64660] = 8'b1110100;
DRAM[64661] = 8'b1110001;
DRAM[64662] = 8'b1111010;
DRAM[64663] = 8'b1101010;
DRAM[64664] = 8'b1101101;
DRAM[64665] = 8'b1101001;
DRAM[64666] = 8'b1101101;
DRAM[64667] = 8'b1111001;
DRAM[64668] = 8'b1111101;
DRAM[64669] = 8'b1110111;
DRAM[64670] = 8'b1110101;
DRAM[64671] = 8'b1111010;
DRAM[64672] = 8'b1111000;
DRAM[64673] = 8'b1110100;
DRAM[64674] = 8'b1110001;
DRAM[64675] = 8'b1110010;
DRAM[64676] = 8'b1111000;
DRAM[64677] = 8'b1111101;
DRAM[64678] = 8'b10000000;
DRAM[64679] = 8'b10000000;
DRAM[64680] = 8'b1111110;
DRAM[64681] = 8'b1111100;
DRAM[64682] = 8'b1111011;
DRAM[64683] = 8'b1111101;
DRAM[64684] = 8'b1111111;
DRAM[64685] = 8'b10000000;
DRAM[64686] = 8'b10000000;
DRAM[64687] = 8'b10000000;
DRAM[64688] = 8'b10000001;
DRAM[64689] = 8'b10000100;
DRAM[64690] = 8'b10001000;
DRAM[64691] = 8'b10001011;
DRAM[64692] = 8'b10001110;
DRAM[64693] = 8'b10010100;
DRAM[64694] = 8'b10011011;
DRAM[64695] = 8'b10100001;
DRAM[64696] = 8'b10110001;
DRAM[64697] = 8'b10110011;
DRAM[64698] = 8'b10111010;
DRAM[64699] = 8'b11000101;
DRAM[64700] = 8'b11001110;
DRAM[64701] = 8'b11010100;
DRAM[64702] = 8'b11011100;
DRAM[64703] = 8'b11100100;
DRAM[64704] = 8'b11101000;
DRAM[64705] = 8'b11101000;
DRAM[64706] = 8'b11010001;
DRAM[64707] = 8'b10110001;
DRAM[64708] = 8'b10100001;
DRAM[64709] = 8'b10010101;
DRAM[64710] = 8'b10000111;
DRAM[64711] = 8'b10000011;
DRAM[64712] = 8'b10000001;
DRAM[64713] = 8'b1111011;
DRAM[64714] = 8'b1111000;
DRAM[64715] = 8'b1111000;
DRAM[64716] = 8'b1110101;
DRAM[64717] = 8'b1101110;
DRAM[64718] = 8'b1101010;
DRAM[64719] = 8'b1101001;
DRAM[64720] = 8'b1100011;
DRAM[64721] = 8'b1100001;
DRAM[64722] = 8'b1011111;
DRAM[64723] = 8'b1011101;
DRAM[64724] = 8'b1011011;
DRAM[64725] = 8'b1011010;
DRAM[64726] = 8'b1011010;
DRAM[64727] = 8'b1011001;
DRAM[64728] = 8'b1011010;
DRAM[64729] = 8'b1011010;
DRAM[64730] = 8'b1011011;
DRAM[64731] = 8'b1011100;
DRAM[64732] = 8'b1011101;
DRAM[64733] = 8'b1011111;
DRAM[64734] = 8'b1100001;
DRAM[64735] = 8'b1100010;
DRAM[64736] = 8'b1100001;
DRAM[64737] = 8'b1100010;
DRAM[64738] = 8'b1100011;
DRAM[64739] = 8'b1100100;
DRAM[64740] = 8'b1100101;
DRAM[64741] = 8'b1100110;
DRAM[64742] = 8'b1100101;
DRAM[64743] = 8'b1100101;
DRAM[64744] = 8'b1100110;
DRAM[64745] = 8'b1100110;
DRAM[64746] = 8'b1100110;
DRAM[64747] = 8'b1100111;
DRAM[64748] = 8'b1100111;
DRAM[64749] = 8'b1101000;
DRAM[64750] = 8'b1101000;
DRAM[64751] = 8'b1101000;
DRAM[64752] = 8'b1101001;
DRAM[64753] = 8'b1101010;
DRAM[64754] = 8'b1101011;
DRAM[64755] = 8'b1101011;
DRAM[64756] = 8'b1101100;
DRAM[64757] = 8'b1101100;
DRAM[64758] = 8'b1101011;
DRAM[64759] = 8'b1101011;
DRAM[64760] = 8'b1101100;
DRAM[64761] = 8'b1101100;
DRAM[64762] = 8'b1101011;
DRAM[64763] = 8'b1101010;
DRAM[64764] = 8'b1101000;
DRAM[64765] = 8'b1100111;
DRAM[64766] = 8'b1100110;
DRAM[64767] = 8'b1100110;
DRAM[64768] = 8'b10001111;
DRAM[64769] = 8'b10001111;
DRAM[64770] = 8'b10010000;
DRAM[64771] = 8'b10010100;
DRAM[64772] = 8'b10011111;
DRAM[64773] = 8'b10110010;
DRAM[64774] = 8'b11001010;
DRAM[64775] = 8'b11011010;
DRAM[64776] = 8'b11101001;
DRAM[64777] = 8'b11101010;
DRAM[64778] = 8'b11101001;
DRAM[64779] = 8'b11101000;
DRAM[64780] = 8'b11100101;
DRAM[64781] = 8'b11100011;
DRAM[64782] = 8'b11100000;
DRAM[64783] = 8'b11011110;
DRAM[64784] = 8'b11100000;
DRAM[64785] = 8'b11100001;
DRAM[64786] = 8'b11100011;
DRAM[64787] = 8'b11100100;
DRAM[64788] = 8'b11100100;
DRAM[64789] = 8'b11011111;
DRAM[64790] = 8'b11010111;
DRAM[64791] = 8'b11010001;
DRAM[64792] = 8'b11001110;
DRAM[64793] = 8'b11001100;
DRAM[64794] = 8'b11001011;
DRAM[64795] = 8'b11001010;
DRAM[64796] = 8'b11001000;
DRAM[64797] = 8'b11000101;
DRAM[64798] = 8'b11000001;
DRAM[64799] = 8'b10111101;
DRAM[64800] = 8'b10111010;
DRAM[64801] = 8'b10111010;
DRAM[64802] = 8'b10111010;
DRAM[64803] = 8'b10111100;
DRAM[64804] = 8'b11000000;
DRAM[64805] = 8'b10111110;
DRAM[64806] = 8'b10110001;
DRAM[64807] = 8'b10100001;
DRAM[64808] = 8'b10101001;
DRAM[64809] = 8'b10101000;
DRAM[64810] = 8'b10100100;
DRAM[64811] = 8'b10011111;
DRAM[64812] = 8'b10011100;
DRAM[64813] = 8'b10011100;
DRAM[64814] = 8'b10011000;
DRAM[64815] = 8'b10010011;
DRAM[64816] = 8'b10010010;
DRAM[64817] = 8'b10010100;
DRAM[64818] = 8'b10010101;
DRAM[64819] = 8'b10010110;
DRAM[64820] = 8'b10010101;
DRAM[64821] = 8'b10010010;
DRAM[64822] = 8'b10001110;
DRAM[64823] = 8'b10001100;
DRAM[64824] = 8'b10010011;
DRAM[64825] = 8'b10010111;
DRAM[64826] = 8'b10011100;
DRAM[64827] = 8'b10011010;
DRAM[64828] = 8'b10010100;
DRAM[64829] = 8'b10001110;
DRAM[64830] = 8'b10001100;
DRAM[64831] = 8'b10001101;
DRAM[64832] = 8'b10001111;
DRAM[64833] = 8'b10001001;
DRAM[64834] = 8'b10001000;
DRAM[64835] = 8'b10001100;
DRAM[64836] = 8'b10001001;
DRAM[64837] = 8'b10000000;
DRAM[64838] = 8'b1111100;
DRAM[64839] = 8'b1111111;
DRAM[64840] = 8'b1111101;
DRAM[64841] = 8'b1111001;
DRAM[64842] = 8'b1110010;
DRAM[64843] = 8'b1101011;
DRAM[64844] = 8'b1100101;
DRAM[64845] = 8'b1100010;
DRAM[64846] = 8'b1100001;
DRAM[64847] = 8'b1100001;
DRAM[64848] = 8'b1101111;
DRAM[64849] = 8'b1011111;
DRAM[64850] = 8'b1010000;
DRAM[64851] = 8'b1010000;
DRAM[64852] = 8'b1011001;
DRAM[64853] = 8'b1100001;
DRAM[64854] = 8'b1100110;
DRAM[64855] = 8'b1101001;
DRAM[64856] = 8'b1111011;
DRAM[64857] = 8'b1101111;
DRAM[64858] = 8'b1110011;
DRAM[64859] = 8'b1101101;
DRAM[64860] = 8'b1101100;
DRAM[64861] = 8'b1101111;
DRAM[64862] = 8'b1100101;
DRAM[64863] = 8'b1101011;
DRAM[64864] = 8'b1110111;
DRAM[64865] = 8'b1101010;
DRAM[64866] = 8'b1100011;
DRAM[64867] = 8'b1101011;
DRAM[64868] = 8'b1110111;
DRAM[64869] = 8'b1111001;
DRAM[64870] = 8'b1110100;
DRAM[64871] = 8'b1101111;
DRAM[64872] = 8'b1101101;
DRAM[64873] = 8'b1110010;
DRAM[64874] = 8'b1110001;
DRAM[64875] = 8'b1101011;
DRAM[64876] = 8'b1101100;
DRAM[64877] = 8'b1110010;
DRAM[64878] = 8'b1101111;
DRAM[64879] = 8'b1101000;
DRAM[64880] = 8'b1101110;
DRAM[64881] = 8'b1101001;
DRAM[64882] = 8'b1100100;
DRAM[64883] = 8'b1100100;
DRAM[64884] = 8'b1100110;
DRAM[64885] = 8'b1100101;
DRAM[64886] = 8'b1100000;
DRAM[64887] = 8'b1011010;
DRAM[64888] = 8'b1100100;
DRAM[64889] = 8'b1100101;
DRAM[64890] = 8'b1100110;
DRAM[64891] = 8'b1100111;
DRAM[64892] = 8'b1101001;
DRAM[64893] = 8'b1101101;
DRAM[64894] = 8'b1110010;
DRAM[64895] = 8'b1110110;
DRAM[64896] = 8'b1111100;
DRAM[64897] = 8'b1101110;
DRAM[64898] = 8'b1100100;
DRAM[64899] = 8'b1100110;
DRAM[64900] = 8'b1100111;
DRAM[64901] = 8'b1100100;
DRAM[64902] = 8'b1101011;
DRAM[64903] = 8'b1111011;
DRAM[64904] = 8'b1100101;
DRAM[64905] = 8'b1100001;
DRAM[64906] = 8'b1101011;
DRAM[64907] = 8'b1110100;
DRAM[64908] = 8'b1110001;
DRAM[64909] = 8'b1110000;
DRAM[64910] = 8'b1110001;
DRAM[64911] = 8'b1101100;
DRAM[64912] = 8'b1110011;
DRAM[64913] = 8'b1110001;
DRAM[64914] = 8'b1101100;
DRAM[64915] = 8'b1111000;
DRAM[64916] = 8'b1110110;
DRAM[64917] = 8'b1110001;
DRAM[64918] = 8'b1111000;
DRAM[64919] = 8'b1100110;
DRAM[64920] = 8'b1110000;
DRAM[64921] = 8'b1101100;
DRAM[64922] = 8'b1101100;
DRAM[64923] = 8'b1110011;
DRAM[64924] = 8'b1110111;
DRAM[64925] = 8'b1110111;
DRAM[64926] = 8'b1110101;
DRAM[64927] = 8'b1110100;
DRAM[64928] = 8'b1111001;
DRAM[64929] = 8'b1110101;
DRAM[64930] = 8'b1110001;
DRAM[64931] = 8'b1110000;
DRAM[64932] = 8'b1110010;
DRAM[64933] = 8'b1110111;
DRAM[64934] = 8'b1111011;
DRAM[64935] = 8'b1111110;
DRAM[64936] = 8'b10000000;
DRAM[64937] = 8'b1111011;
DRAM[64938] = 8'b1111001;
DRAM[64939] = 8'b1111100;
DRAM[64940] = 8'b1111110;
DRAM[64941] = 8'b1111110;
DRAM[64942] = 8'b1111111;
DRAM[64943] = 8'b10000001;
DRAM[64944] = 8'b10000011;
DRAM[64945] = 8'b10000110;
DRAM[64946] = 8'b10001011;
DRAM[64947] = 8'b10001110;
DRAM[64948] = 8'b10010010;
DRAM[64949] = 8'b10010110;
DRAM[64950] = 8'b10011011;
DRAM[64951] = 8'b10011111;
DRAM[64952] = 8'b10101100;
DRAM[64953] = 8'b10101100;
DRAM[64954] = 8'b10110011;
DRAM[64955] = 8'b10111111;
DRAM[64956] = 8'b11001010;
DRAM[64957] = 8'b11010001;
DRAM[64958] = 8'b11011001;
DRAM[64959] = 8'b11100000;
DRAM[64960] = 8'b11100110;
DRAM[64961] = 8'b11101001;
DRAM[64962] = 8'b11011001;
DRAM[64963] = 8'b11000010;
DRAM[64964] = 8'b10110111;
DRAM[64965] = 8'b10101000;
DRAM[64966] = 8'b10010010;
DRAM[64967] = 8'b10000110;
DRAM[64968] = 8'b10001010;
DRAM[64969] = 8'b10000010;
DRAM[64970] = 8'b1111011;
DRAM[64971] = 8'b1111000;
DRAM[64972] = 8'b1110010;
DRAM[64973] = 8'b1101010;
DRAM[64974] = 8'b1100101;
DRAM[64975] = 8'b1100100;
DRAM[64976] = 8'b1100010;
DRAM[64977] = 8'b1100001;
DRAM[64978] = 8'b1011110;
DRAM[64979] = 8'b1011100;
DRAM[64980] = 8'b1011010;
DRAM[64981] = 8'b1011000;
DRAM[64982] = 8'b1010111;
DRAM[64983] = 8'b1010111;
DRAM[64984] = 8'b1011010;
DRAM[64985] = 8'b1011010;
DRAM[64986] = 8'b1011010;
DRAM[64987] = 8'b1011011;
DRAM[64988] = 8'b1011101;
DRAM[64989] = 8'b1011111;
DRAM[64990] = 8'b1100001;
DRAM[64991] = 8'b1100010;
DRAM[64992] = 8'b1100001;
DRAM[64993] = 8'b1100010;
DRAM[64994] = 8'b1100011;
DRAM[64995] = 8'b1100100;
DRAM[64996] = 8'b1100101;
DRAM[64997] = 8'b1100110;
DRAM[64998] = 8'b1100101;
DRAM[64999] = 8'b1100101;
DRAM[65000] = 8'b1100110;
DRAM[65001] = 8'b1100110;
DRAM[65002] = 8'b1100110;
DRAM[65003] = 8'b1100111;
DRAM[65004] = 8'b1100111;
DRAM[65005] = 8'b1101000;
DRAM[65006] = 8'b1101000;
DRAM[65007] = 8'b1101000;
DRAM[65008] = 8'b1101001;
DRAM[65009] = 8'b1101001;
DRAM[65010] = 8'b1101010;
DRAM[65011] = 8'b1101011;
DRAM[65012] = 8'b1101011;
DRAM[65013] = 8'b1101011;
DRAM[65014] = 8'b1101011;
DRAM[65015] = 8'b1101011;
DRAM[65016] = 8'b1101100;
DRAM[65017] = 8'b1101100;
DRAM[65018] = 8'b1101011;
DRAM[65019] = 8'b1101010;
DRAM[65020] = 8'b1101000;
DRAM[65021] = 8'b1100111;
DRAM[65022] = 8'b1100110;
DRAM[65023] = 8'b1100110;
DRAM[65024] = 8'b10001101;
DRAM[65025] = 8'b10010000;
DRAM[65026] = 8'b10010101;
DRAM[65027] = 8'b10011011;
DRAM[65028] = 8'b10101000;
DRAM[65029] = 8'b10111101;
DRAM[65030] = 8'b11010010;
DRAM[65031] = 8'b11100000;
DRAM[65032] = 8'b11101001;
DRAM[65033] = 8'b11100110;
DRAM[65034] = 8'b11100101;
DRAM[65035] = 8'b11100100;
DRAM[65036] = 8'b11100011;
DRAM[65037] = 8'b11100000;
DRAM[65038] = 8'b11011110;
DRAM[65039] = 8'b11011110;
DRAM[65040] = 8'b11011110;
DRAM[65041] = 8'b11011111;
DRAM[65042] = 8'b11100000;
DRAM[65043] = 8'b11100010;
DRAM[65044] = 8'b11100001;
DRAM[65045] = 8'b11011100;
DRAM[65046] = 8'b11010100;
DRAM[65047] = 8'b11001111;
DRAM[65048] = 8'b11001101;
DRAM[65049] = 8'b11001011;
DRAM[65050] = 8'b11001010;
DRAM[65051] = 8'b11001001;
DRAM[65052] = 8'b11001000;
DRAM[65053] = 8'b11000100;
DRAM[65054] = 8'b11000000;
DRAM[65055] = 8'b10111100;
DRAM[65056] = 8'b10111101;
DRAM[65057] = 8'b11000000;
DRAM[65058] = 8'b11000001;
DRAM[65059] = 8'b10111100;
DRAM[65060] = 8'b10110111;
DRAM[65061] = 8'b10110001;
DRAM[65062] = 8'b10101000;
DRAM[65063] = 8'b10011111;
DRAM[65064] = 8'b10100001;
DRAM[65065] = 8'b10100001;
DRAM[65066] = 8'b10011100;
DRAM[65067] = 8'b10010101;
DRAM[65068] = 8'b10010011;
DRAM[65069] = 8'b10010101;
DRAM[65070] = 8'b10010011;
DRAM[65071] = 8'b10001110;
DRAM[65072] = 8'b10001111;
DRAM[65073] = 8'b10001110;
DRAM[65074] = 8'b10001101;
DRAM[65075] = 8'b10001100;
DRAM[65076] = 8'b10001101;
DRAM[65077] = 8'b10001111;
DRAM[65078] = 8'b10010001;
DRAM[65079] = 8'b10010011;
DRAM[65080] = 8'b10011101;
DRAM[65081] = 8'b10011000;
DRAM[65082] = 8'b10010010;
DRAM[65083] = 8'b10001110;
DRAM[65084] = 8'b10001100;
DRAM[65085] = 8'b10001011;
DRAM[65086] = 8'b10001001;
DRAM[65087] = 8'b10000111;
DRAM[65088] = 8'b10001111;
DRAM[65089] = 8'b10001010;
DRAM[65090] = 8'b10000111;
DRAM[65091] = 8'b10000110;
DRAM[65092] = 8'b10000011;
DRAM[65093] = 8'b1111100;
DRAM[65094] = 8'b1110011;
DRAM[65095] = 8'b1101110;
DRAM[65096] = 8'b1101000;
DRAM[65097] = 8'b1101100;
DRAM[65098] = 8'b1110001;
DRAM[65099] = 8'b1110011;
DRAM[65100] = 8'b1101111;
DRAM[65101] = 8'b1100110;
DRAM[65102] = 8'b1011011;
DRAM[65103] = 8'b1010100;
DRAM[65104] = 8'b1110010;
DRAM[65105] = 8'b1101001;
DRAM[65106] = 8'b1011010;
DRAM[65107] = 8'b1001110;
DRAM[65108] = 8'b1001110;
DRAM[65109] = 8'b1011011;
DRAM[65110] = 8'b1101000;
DRAM[65111] = 8'b1101110;
DRAM[65112] = 8'b1111000;
DRAM[65113] = 8'b1101011;
DRAM[65114] = 8'b1110000;
DRAM[65115] = 8'b1101111;
DRAM[65116] = 8'b1110001;
DRAM[65117] = 8'b1110001;
DRAM[65118] = 8'b1100010;
DRAM[65119] = 8'b1100110;
DRAM[65120] = 8'b1110100;
DRAM[65121] = 8'b1101100;
DRAM[65122] = 8'b1100111;
DRAM[65123] = 8'b1101001;
DRAM[65124] = 8'b1101110;
DRAM[65125] = 8'b1110000;
DRAM[65126] = 8'b1110000;
DRAM[65127] = 8'b1110000;
DRAM[65128] = 8'b1101011;
DRAM[65129] = 8'b1101101;
DRAM[65130] = 8'b1101111;
DRAM[65131] = 8'b1101100;
DRAM[65132] = 8'b1100111;
DRAM[65133] = 8'b1100100;
DRAM[65134] = 8'b1101000;
DRAM[65135] = 8'b1101101;
DRAM[65136] = 8'b1101011;
DRAM[65137] = 8'b1100101;
DRAM[65138] = 8'b1100001;
DRAM[65139] = 8'b1100100;
DRAM[65140] = 8'b1101011;
DRAM[65141] = 8'b1101101;
DRAM[65142] = 8'b1101001;
DRAM[65143] = 8'b1100011;
DRAM[65144] = 8'b1100100;
DRAM[65145] = 8'b1100100;
DRAM[65146] = 8'b1100100;
DRAM[65147] = 8'b1101000;
DRAM[65148] = 8'b1101101;
DRAM[65149] = 8'b1110010;
DRAM[65150] = 8'b1110101;
DRAM[65151] = 8'b1110110;
DRAM[65152] = 8'b1111001;
DRAM[65153] = 8'b1110110;
DRAM[65154] = 8'b1101000;
DRAM[65155] = 8'b1100110;
DRAM[65156] = 8'b1101110;
DRAM[65157] = 8'b1100101;
DRAM[65158] = 8'b1100011;
DRAM[65159] = 8'b1111010;
DRAM[65160] = 8'b1101010;
DRAM[65161] = 8'b1100001;
DRAM[65162] = 8'b1101000;
DRAM[65163] = 8'b1110101;
DRAM[65164] = 8'b1110101;
DRAM[65165] = 8'b1110100;
DRAM[65166] = 8'b1110010;
DRAM[65167] = 8'b1101010;
DRAM[65168] = 8'b1110010;
DRAM[65169] = 8'b1110001;
DRAM[65170] = 8'b1101100;
DRAM[65171] = 8'b1111001;
DRAM[65172] = 8'b1111000;
DRAM[65173] = 8'b1110011;
DRAM[65174] = 8'b1110111;
DRAM[65175] = 8'b1100100;
DRAM[65176] = 8'b1101100;
DRAM[65177] = 8'b1101100;
DRAM[65178] = 8'b1101011;
DRAM[65179] = 8'b1101100;
DRAM[65180] = 8'b1110010;
DRAM[65181] = 8'b1110111;
DRAM[65182] = 8'b1110100;
DRAM[65183] = 8'b1101100;
DRAM[65184] = 8'b1110111;
DRAM[65185] = 8'b1110101;
DRAM[65186] = 8'b1110000;
DRAM[65187] = 8'b1101100;
DRAM[65188] = 8'b1101100;
DRAM[65189] = 8'b1101111;
DRAM[65190] = 8'b1110110;
DRAM[65191] = 8'b1111011;
DRAM[65192] = 8'b10000000;
DRAM[65193] = 8'b1111010;
DRAM[65194] = 8'b1110111;
DRAM[65195] = 8'b1111100;
DRAM[65196] = 8'b1111111;
DRAM[65197] = 8'b1111111;
DRAM[65198] = 8'b10000001;
DRAM[65199] = 8'b10000110;
DRAM[65200] = 8'b10000101;
DRAM[65201] = 8'b10001000;
DRAM[65202] = 8'b10001101;
DRAM[65203] = 8'b10010010;
DRAM[65204] = 8'b10010110;
DRAM[65205] = 8'b10011001;
DRAM[65206] = 8'b10011100;
DRAM[65207] = 8'b10011110;
DRAM[65208] = 8'b10100101;
DRAM[65209] = 8'b10100100;
DRAM[65210] = 8'b10101001;
DRAM[65211] = 8'b10110101;
DRAM[65212] = 8'b11000000;
DRAM[65213] = 8'b11001000;
DRAM[65214] = 8'b11010001;
DRAM[65215] = 8'b11011000;
DRAM[65216] = 8'b11100110;
DRAM[65217] = 8'b11100110;
DRAM[65218] = 8'b11010001;
DRAM[65219] = 8'b10110110;
DRAM[65220] = 8'b10101100;
DRAM[65221] = 8'b10100011;
DRAM[65222] = 8'b10010100;
DRAM[65223] = 8'b10001101;
DRAM[65224] = 8'b10001011;
DRAM[65225] = 8'b10000011;
DRAM[65226] = 8'b1111010;
DRAM[65227] = 8'b1110101;
DRAM[65228] = 8'b1110000;
DRAM[65229] = 8'b1101000;
DRAM[65230] = 8'b1100101;
DRAM[65231] = 8'b1100101;
DRAM[65232] = 8'b1100010;
DRAM[65233] = 8'b1100001;
DRAM[65234] = 8'b1011110;
DRAM[65235] = 8'b1011011;
DRAM[65236] = 8'b1011000;
DRAM[65237] = 8'b1010110;
DRAM[65238] = 8'b1010101;
DRAM[65239] = 8'b1010100;
DRAM[65240] = 8'b1011000;
DRAM[65241] = 8'b1011000;
DRAM[65242] = 8'b1011001;
DRAM[65243] = 8'b1011010;
DRAM[65244] = 8'b1011011;
DRAM[65245] = 8'b1011101;
DRAM[65246] = 8'b1011111;
DRAM[65247] = 8'b1100000;
DRAM[65248] = 8'b1100001;
DRAM[65249] = 8'b1100010;
DRAM[65250] = 8'b1100011;
DRAM[65251] = 8'b1100100;
DRAM[65252] = 8'b1100101;
DRAM[65253] = 8'b1100110;
DRAM[65254] = 8'b1100101;
DRAM[65255] = 8'b1100101;
DRAM[65256] = 8'b1100110;
DRAM[65257] = 8'b1100110;
DRAM[65258] = 8'b1100110;
DRAM[65259] = 8'b1100111;
DRAM[65260] = 8'b1100111;
DRAM[65261] = 8'b1101000;
DRAM[65262] = 8'b1101000;
DRAM[65263] = 8'b1101000;
DRAM[65264] = 8'b1101000;
DRAM[65265] = 8'b1101001;
DRAM[65266] = 8'b1101010;
DRAM[65267] = 8'b1101011;
DRAM[65268] = 8'b1101011;
DRAM[65269] = 8'b1101011;
DRAM[65270] = 8'b1101011;
DRAM[65271] = 8'b1101010;
DRAM[65272] = 8'b1101100;
DRAM[65273] = 8'b1101100;
DRAM[65274] = 8'b1101011;
DRAM[65275] = 8'b1101010;
DRAM[65276] = 8'b1101000;
DRAM[65277] = 8'b1100111;
DRAM[65278] = 8'b1100110;
DRAM[65279] = 8'b1100110;
DRAM[65280] = 8'b10001111;
DRAM[65281] = 8'b10010100;
DRAM[65282] = 8'b10011010;
DRAM[65283] = 8'b10100011;
DRAM[65284] = 8'b10110001;
DRAM[65285] = 8'b11000110;
DRAM[65286] = 8'b11011010;
DRAM[65287] = 8'b11100101;
DRAM[65288] = 8'b11100111;
DRAM[65289] = 8'b11100100;
DRAM[65290] = 8'b11100001;
DRAM[65291] = 8'b11100001;
DRAM[65292] = 8'b11100001;
DRAM[65293] = 8'b11011110;
DRAM[65294] = 8'b11011101;
DRAM[65295] = 8'b11011101;
DRAM[65296] = 8'b11011100;
DRAM[65297] = 8'b11011101;
DRAM[65298] = 8'b11011111;
DRAM[65299] = 8'b11100000;
DRAM[65300] = 8'b11011111;
DRAM[65301] = 8'b11011010;
DRAM[65302] = 8'b11010010;
DRAM[65303] = 8'b11001100;
DRAM[65304] = 8'b11001001;
DRAM[65305] = 8'b11000111;
DRAM[65306] = 8'b11000110;
DRAM[65307] = 8'b11000110;
DRAM[65308] = 8'b11000100;
DRAM[65309] = 8'b11000001;
DRAM[65310] = 8'b10111100;
DRAM[65311] = 8'b10111000;
DRAM[65312] = 8'b10101110;
DRAM[65313] = 8'b10111000;
DRAM[65314] = 8'b10111101;
DRAM[65315] = 8'b10110111;
DRAM[65316] = 8'b10101110;
DRAM[65317] = 8'b10101011;
DRAM[65318] = 8'b10101100;
DRAM[65319] = 8'b10101100;
DRAM[65320] = 8'b10011011;
DRAM[65321] = 8'b10011010;
DRAM[65322] = 8'b10010101;
DRAM[65323] = 8'b10001101;
DRAM[65324] = 8'b10001101;
DRAM[65325] = 8'b10010011;
DRAM[65326] = 8'b10010101;
DRAM[65327] = 8'b10010001;
DRAM[65328] = 8'b10001010;
DRAM[65329] = 8'b10000111;
DRAM[65330] = 8'b10000010;
DRAM[65331] = 8'b1111111;
DRAM[65332] = 8'b10000000;
DRAM[65333] = 8'b10000110;
DRAM[65334] = 8'b10001100;
DRAM[65335] = 8'b10010001;
DRAM[65336] = 8'b10011001;
DRAM[65337] = 8'b10001101;
DRAM[65338] = 8'b10000001;
DRAM[65339] = 8'b10000000;
DRAM[65340] = 8'b10001001;
DRAM[65341] = 8'b10010010;
DRAM[65342] = 8'b10010011;
DRAM[65343] = 8'b10010001;
DRAM[65344] = 8'b10001000;
DRAM[65345] = 8'b10000011;
DRAM[65346] = 8'b1111101;
DRAM[65347] = 8'b1111001;
DRAM[65348] = 8'b1111100;
DRAM[65349] = 8'b1111111;
DRAM[65350] = 8'b1111101;
DRAM[65351] = 8'b1110111;
DRAM[65352] = 8'b1101000;
DRAM[65353] = 8'b1101010;
DRAM[65354] = 8'b1101110;
DRAM[65355] = 8'b1110000;
DRAM[65356] = 8'b1101111;
DRAM[65357] = 8'b1101101;
DRAM[65358] = 8'b1101001;
DRAM[65359] = 8'b1100110;
DRAM[65360] = 8'b1000110;
DRAM[65361] = 8'b1100000;
DRAM[65362] = 8'b1110000;
DRAM[65363] = 8'b1101001;
DRAM[65364] = 8'b1011100;
DRAM[65365] = 8'b1011101;
DRAM[65366] = 8'b1101000;
DRAM[65367] = 8'b1101111;
DRAM[65368] = 8'b1110111;
DRAM[65369] = 8'b1101000;
DRAM[65370] = 8'b1101110;
DRAM[65371] = 8'b1101111;
DRAM[65372] = 8'b1110100;
DRAM[65373] = 8'b1110011;
DRAM[65374] = 8'b1100001;
DRAM[65375] = 8'b1100011;
DRAM[65376] = 8'b1101111;
DRAM[65377] = 8'b1101101;
DRAM[65378] = 8'b1101011;
DRAM[65379] = 8'b1101010;
DRAM[65380] = 8'b1101000;
DRAM[65381] = 8'b1100110;
DRAM[65382] = 8'b1101010;
DRAM[65383] = 8'b1101110;
DRAM[65384] = 8'b1111000;
DRAM[65385] = 8'b1101011;
DRAM[65386] = 8'b1101000;
DRAM[65387] = 8'b1110000;
DRAM[65388] = 8'b1110000;
DRAM[65389] = 8'b1100110;
DRAM[65390] = 8'b1100110;
DRAM[65391] = 8'b1110010;
DRAM[65392] = 8'b1101001;
DRAM[65393] = 8'b1100011;
DRAM[65394] = 8'b1011110;
DRAM[65395] = 8'b1100000;
DRAM[65396] = 8'b1100111;
DRAM[65397] = 8'b1101010;
DRAM[65398] = 8'b1100111;
DRAM[65399] = 8'b1100011;
DRAM[65400] = 8'b1101011;
DRAM[65401] = 8'b1101000;
DRAM[65402] = 8'b1100110;
DRAM[65403] = 8'b1101000;
DRAM[65404] = 8'b1101101;
DRAM[65405] = 8'b1101111;
DRAM[65406] = 8'b1101111;
DRAM[65407] = 8'b1101101;
DRAM[65408] = 8'b1110011;
DRAM[65409] = 8'b1111101;
DRAM[65410] = 8'b1101011;
DRAM[65411] = 8'b1100010;
DRAM[65412] = 8'b1101110;
DRAM[65413] = 8'b1100011;
DRAM[65414] = 8'b1011001;
DRAM[65415] = 8'b1101110;
DRAM[65416] = 8'b1101111;
DRAM[65417] = 8'b1100010;
DRAM[65418] = 8'b1100111;
DRAM[65419] = 8'b1110101;
DRAM[65420] = 8'b1111000;
DRAM[65421] = 8'b1110111;
DRAM[65422] = 8'b1110011;
DRAM[65423] = 8'b1101001;
DRAM[65424] = 8'b1110000;
DRAM[65425] = 8'b1101111;
DRAM[65426] = 8'b1101100;
DRAM[65427] = 8'b1111010;
DRAM[65428] = 8'b1111010;
DRAM[65429] = 8'b1110101;
DRAM[65430] = 8'b1111000;
DRAM[65431] = 8'b1100011;
DRAM[65432] = 8'b1100111;
DRAM[65433] = 8'b1101011;
DRAM[65434] = 8'b1101010;
DRAM[65435] = 8'b1101001;
DRAM[65436] = 8'b1110000;
DRAM[65437] = 8'b1111000;
DRAM[65438] = 8'b1110011;
DRAM[65439] = 8'b1100110;
DRAM[65440] = 8'b1110101;
DRAM[65441] = 8'b1110100;
DRAM[65442] = 8'b1110000;
DRAM[65443] = 8'b1101010;
DRAM[65444] = 8'b1100111;
DRAM[65445] = 8'b1101001;
DRAM[65446] = 8'b1110001;
DRAM[65447] = 8'b1111000;
DRAM[65448] = 8'b1111000;
DRAM[65449] = 8'b1110001;
DRAM[65450] = 8'b1101111;
DRAM[65451] = 8'b1110101;
DRAM[65452] = 8'b1111010;
DRAM[65453] = 8'b1111010;
DRAM[65454] = 8'b1111110;
DRAM[65455] = 8'b10000100;
DRAM[65456] = 8'b10000000;
DRAM[65457] = 8'b10000100;
DRAM[65458] = 8'b10001001;
DRAM[65459] = 8'b10001111;
DRAM[65460] = 8'b10010100;
DRAM[65461] = 8'b10010110;
DRAM[65462] = 8'b10011000;
DRAM[65463] = 8'b10011001;
DRAM[65464] = 8'b10100101;
DRAM[65465] = 8'b10100011;
DRAM[65466] = 8'b10100111;
DRAM[65467] = 8'b10110011;
DRAM[65468] = 8'b10111110;
DRAM[65469] = 8'b11000110;
DRAM[65470] = 8'b11001111;
DRAM[65471] = 8'b11010110;
DRAM[65472] = 8'b11100111;
DRAM[65473] = 8'b11100001;
DRAM[65474] = 8'b11000000;
DRAM[65475] = 8'b10011100;
DRAM[65476] = 8'b10010000;
DRAM[65477] = 8'b10001111;
DRAM[65478] = 8'b10001111;
DRAM[65479] = 8'b10010011;
DRAM[65480] = 8'b10000111;
DRAM[65481] = 8'b1111110;
DRAM[65482] = 8'b1110110;
DRAM[65483] = 8'b1110010;
DRAM[65484] = 8'b1101111;
DRAM[65485] = 8'b1101010;
DRAM[65486] = 8'b1101000;
DRAM[65487] = 8'b1101010;
DRAM[65488] = 8'b1100011;
DRAM[65489] = 8'b1100001;
DRAM[65490] = 8'b1011110;
DRAM[65491] = 8'b1011011;
DRAM[65492] = 8'b1010111;
DRAM[65493] = 8'b1010101;
DRAM[65494] = 8'b1010100;
DRAM[65495] = 8'b1010011;
DRAM[65496] = 8'b1010111;
DRAM[65497] = 8'b1010111;
DRAM[65498] = 8'b1010111;
DRAM[65499] = 8'b1011000;
DRAM[65500] = 8'b1011010;
DRAM[65501] = 8'b1011100;
DRAM[65502] = 8'b1011110;
DRAM[65503] = 8'b1011111;
DRAM[65504] = 8'b1100001;
DRAM[65505] = 8'b1100010;
DRAM[65506] = 8'b1100011;
DRAM[65507] = 8'b1100100;
DRAM[65508] = 8'b1100101;
DRAM[65509] = 8'b1100110;
DRAM[65510] = 8'b1100101;
DRAM[65511] = 8'b1100101;
DRAM[65512] = 8'b1100110;
DRAM[65513] = 8'b1100110;
DRAM[65514] = 8'b1100110;
DRAM[65515] = 8'b1100111;
DRAM[65516] = 8'b1100111;
DRAM[65517] = 8'b1101000;
DRAM[65518] = 8'b1101000;
DRAM[65519] = 8'b1101000;
DRAM[65520] = 8'b1101000;
DRAM[65521] = 8'b1101001;
DRAM[65522] = 8'b1101010;
DRAM[65523] = 8'b1101011;
DRAM[65524] = 8'b1101011;
DRAM[65525] = 8'b1101011;
DRAM[65526] = 8'b1101011;
DRAM[65527] = 8'b1101010;
DRAM[65528] = 8'b1101100;
DRAM[65529] = 8'b1101100;
DRAM[65530] = 8'b1101011;
DRAM[65531] = 8'b1101010;
DRAM[65532] = 8'b1101000;
DRAM[65533] = 8'b1100111;
DRAM[65534] = 8'b1100110;
DRAM[65535] = 8'b1100110;
end

always @ (negedge clock)
begin
    if(wren == 0)
        q <= DRAM[address];
    else
        DRAM[address] <= data;
end
endmodule